library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity TPG is
	generic	(
			 PixelNumber		: std_logic_vector(31 downto 0) := x"00000000"
			 -- Row				: std_logic_vector(11 downto 0) := x"000";
			 -- Column				: std_logic_vector(11 downto 0) := x"000"
			);
	port(
		 nReset   				: in std_logic;
		 Clk     				: in std_logic;
--*********************** Global signals *****************************************
		 s0_read				: in std_logic;
		 -- s0_write				: in std_logic;
		 s0_chipselect			: in std_logic;
		 s0_address				: in std_logic_vector(1 downto 0);
		 s0_readdata			: buffer std_logic_vector(15 downto 0);
		 -- s0_readdatavalid		: out std_logic;
		 -- s0_writedata			: in std_logic_vector(15 downto 0);
		 -- s0_waitrequest			: out std_logic;
--************************* Avalon-MM Slave **************************************
		 Int     				: buffer std_logic--;--interrupt on VSync
--*********************** External signals ***************************************
		);
end TPG;

ARCHITECTURE Arc_TPG OF TPG IS

	-- subtype Video4xPixel is std_logic_vector(31 downto 0);
	-- type Video is array (0 to 76799) of Video4xPixel;
	
	-- signal	VideoData	: Video :=	(
									 -- x"9E9C9A9E", x"A3A19DA0", x"9EA1A5AA", x"AEAFAEAD", x"ACAAAAAD", x"AFAFAEAE", x"B1B1B0AF", x"AFAFAFAF",
									 -- x"AEAFAFB0", x"B3B6B3AF", x"B2B3B4B6", x"B8B9BABB", x"BDBDBDBF", x"C1C3C4C3", x"C4C4C5C5", x"C5C5C4C4",
									 -- x"C5C7C9C9", x"C8C7C8C8", x"C7C8C9C7", x"C6C6C5C3", x"C4C4C3C3", x"C3C4C4C5", x"C4C3C2C1", x"C0BFBEBD",
									 -- x"C0C0C1C1", x"C1C1C0C0", x"C1C1C2C2", x"C2C2C3C4", x"C6C2C4C9", x"CBC8CACF", x"C8C9C9C9", x"C7C7C8C9",
									 -- x"C7C9CCCE", x"CDCDCDCE", x"CFCFCFCD", x"CCCBCBCC", x"C8C9C7C5", x"C5C7C7C5", x"C5C4C4C4", x"C3C2C3C6",
									 -- x"C2C4C4C2", x"C1C1C0BD", x"C1BEBEBF", x"C0BEBEBF", x"C1C2C2C2", x"C2C2C3C4", x"C1C2C3C4", x"C5C6C7C7",
									 -- x"C4CACCCB", x"CACCCCC9", x"CDCAC8C9", x"C9C9CCD0", x"C9CCCECD", x"CBCBCAC9", x"C9C7C6C6", x"C4C1C1C2",
									 -- x"C3C3C4C4", x"C3C2C2C1", x"C3C2C1BF", x"BEBDBDBD", x"BDBEBEBE", x"BDBEBEBF", x"C0C2C2BF", x"BEBEBDBB",
									 -- x"BFBFBEBC", x"B8B4B3B4", x"B2AFA9A4", x"9F9B9897", x"92909092", x"93908D8C", x"8C8C8B8A", x"8C8D8B87",
									 -- x"87888A8B", x"8B8B8B8B", x"8B8B8B8E", x"9091908E", x"9191908E", x"8D8C8C8D", x"8B8B8783", x"8284817C",
									 -- x"7B7B7B7C", x"7B797A7C", x"7D7D7D7C", x"7A797A7C", x"78797A7B", x"7C7C7D7D", x"7D7D7D7C", x"7B7B7B7C",
									 -- x"7D7B7C7C", x"7B7D7D77", x"7B807E7E", x"7A777D7F", x"7B83807A", x"7D7F818A", x"84828182", x"85868684",
									 -- x"83818889", x"83848987", x"878C8C89", x"898D8D88", x"878C8C87", x"878B8C89", x"8688908A", x"8C958E8C",
									 -- x"8C8C8E90", x"8F8C8D90", x"8F909193", x"928F8D8B", x"938F8987", x"8B8B8A8E", x"8C83848A", x"88898C88",
									 -- x"888A8787", x"85868981", x"83898C8A", x"898B8A86", x"85898B89", x"8A8E8E8B", x"888D8B87", x"8A8E8B88",
									 -- x"8E8C8E8E", x"8C93968F", x"93918F90", x"94929196", x"97979AA0", x"A3A1A2A6", x"A4A7A7A7", x"AAABABAF",
									 -- x"A9A6ABA7", x"A8AEA7A7", x"AAA7ABAD", x"A8ABB1AF", x"ABAFB0AD", x"ADAFAFAB", x"ABAFB2B0", x"ABA9ABAF",
									 -- x"ADB1B1AD", x"ADB1AFAA", x"B0ACAEAE", x"ADB3B6B0", x"B3B1B3B7", x"B6B1B0B3", x"AFAFB2B4", x"B3B0B0B3",
									 -- x"B5B5B5B5", x"B4B4B4B3", x"AFB4B6AF", x"ABB3B8B3", x"B7B5B4B6", x"B6B5B6B9", x"B3B5B6B5", x"B4B4B7BA",
									 -- x"BAB6B8BA", x"BBBDBEBB", x"BDBCBCBC", x"BDBDBDBC", x"BBBABAB9", x"B9B9BABA", x"BAB6B5BA", x"BCB9B6B6",
									 -- x"9B9B999B", x"9F9F9D9F", x"A0A2A5A9", x"ABADACAC", x"ADACACAF", x"B0AFAEAF", x"ACACADAE", x"AFAFAFAF",
									 -- x"AEB0B1B1", x"B2B4B2AF", x"B4B4B4B5", x"B6B8BABB", x"BFBEBEC0", x"C3C5C5C4", x"C3C3C4C5", x"C5C5C5C5",
									 -- x"C6C7C7C7", x"C7C7C7C7", x"C7C8C9C8", x"C7C8C7C5", x"C5C5C5C6", x"C5C5C4C4", x"C5C4C2C0", x"C0C1C1C1",
									 -- x"C0C0C1C1", x"C1C1C1C1", x"C1C1C2C2", x"C2C2C3C4", x"C4C2C4C8", x"C9C7C9CC", x"C9CACAC9", x"C8C7C8C9",
									 -- x"C8C9CBCC", x"CDCECECF", x"CFCFCFCE", x"CCCBCBCC", x"C9CAC8C6", x"C5C7C6C4", x"C6C5C4C4", x"C3C2C3C6",
									 -- x"C4C5C4C1", x"C0C1C0BF", x"C2BFBFC1", x"C1C0C0C2", x"C0C1C1C1", x"C1C1C2C3", x"C2C3C3C4", x"C5C6C6C6",
									 -- x"C5CACCCA", x"CACCCCC9", x"CCC9C8C8", x"C9C9CBCE", x"CCCDCDCC", x"CBCCCAC8", x"C9C7C6C7", x"C6C3C3C4",
									 -- x"C5C4C4C3", x"C3C2C1C0", x"C2C2C1C0", x"BFBEBDBC", x"BDBDBEBE", x"BEBEBFC0", x"C0C2C2BF", x"BDBDBDBC",
									 -- x"BFBEBEBD", x"B9B5B4B6", x"B3B0ACA6", x"A29E9A98", x"96939295", x"95939090", x"8D8D8C8A", x"8A8A8988",
									 -- x"88898B8C", x"8C8C8C8C", x"8C8B8C8E", x"9192918F", x"90908F8E", x"8C8B8C8C", x"88888785", x"84827D78",
									 -- x"7A7B7E81", x"7F7D7D7E", x"80807E7C", x"7A797A7B", x"7B7A7A7B", x"7C7C7B7A", x"7F808180", x"7D7A7979",
									 -- x"7C7B7D7F", x"7F82827D", x"7E828182", x"7F7B7F7E", x"79807E7A", x"7D7E7F86", x"84838283", x"84868787",
									 -- x"87838687", x"83858884", x"878B8A86", x"868A8A86", x"898B8A88", x"8A8D8D8B", x"8A8A918D", x"8E928C8B",
									 -- x"8C8B8C8E", x"8F8E8E8F", x"8F8F8F8F", x"8F8D8A89", x"8E8C8887", x"8A89888C", x"8F88898C", x"8A8B8C87",
									 -- x"88898789", x"87878B84", x"898B8C8D", x"8B898989", x"84858789", x"89878585", x"86878484", x"8A8C8B8C",
									 -- x"8B898A8A", x"8B909290", x"9393908F", x"92919093", x"98989B9F", x"A09EA0A5", x"A9A8A7AA", x"AEAAA8AD",
									 -- x"A5A5ACA8", x"A7AAA5A7", x"A9ACB0AF", x"A9A9AFB3", x"ADB1B2B0", x"AEB0B0AD", x"B0B1B3B2", x"B0AFB0B1",
									 -- x"ACADADAD", x"ADADACAA", x"B1B0B0B0", x"B1B5B6B2", x"B3B2B4B7", x"B5B1B0B2", x"B2B1B1B2", x"B0AEB0B4",
									 -- x"B3B4B4B4", x"B5B5B5B5", x"B4B5B6B3", x"AEB1B5B4", x"B6B5B4B6", x"B6B6B7B9", x"BAB9B8B7", x"B7B8B9BA",
									 -- x"BBB8B9BA", x"BABDBFBC", x"BDBDBDBD", x"BDBCBAB9", x"BBBABABA", x"BBBBBCBC", x"BCB9B8BA", x"BBBAB7B5",
									 -- x"9B9E9C9B", x"9E9F9EA0", x"A1A2A4A6", x"A8AAAAAB", x"AEAEAFB0", x"B0AEAEAF", x"AFAFAFAF", x"AFAFAEAE",
									 -- x"ADB0B3B3", x"B2B2B2B1", x"B5B5B4B5", x"B6B7B9BA", x"BFBEBFC1", x"C3C5C4C4", x"C1C2C4C5", x"C6C6C6C5",
									 -- x"C8C7C6C6", x"C6C7C6C6", x"C5C7C8C7", x"C7C8C8C6", x"C5C5C5C5", x"C5C5C5C5", x"C5C3C1BF", x"C0C1C3C4",
									 -- x"C0C1C1C1", x"C1C1C1C0", x"C0C1C2C2", x"C1C2C2C3", x"C1C3C4C5", x"C6C7C8C8", x"CACACAC9", x"C8C7C7C8",
									 -- x"C9C9C9CB", x"CDCFCFD0", x"CFCFCFCE", x"CDCCCCCC", x"CBCAC9C6", x"C6C6C6C4", x"C8C6C5C4", x"C3C2C3C6",
									 -- x"C4C4C3C1", x"C0C1C1C0", x"C1C0BFC1", x"C2C2C2C3", x"C1C2C2C2", x"C2C3C4C5", x"C3C3C4C4", x"C5C5C5C5",
									 -- x"C6C9CBC9", x"C9CBCBC9", x"CAC8C7C8", x"C8C8C9CB", x"CECDCBC9", x"CACBC8C5", x"C6C5C5C6", x"C6C4C4C4",
									 -- x"C6C5C4C3", x"C2C1C0C0", x"C1C1C1C1", x"C0BFBDBC", x"BEBEBEBE", x"BEBEBFC0", x"C1C2C1BF", x"BDBDBDBC",
									 -- x"BDBCBCBB", x"B8B5B4B6", x"B4B2ADA9", x"A5A19D9B", x"98969596", x"97969594", x"9293918D", x"8B8B8C8B",
									 -- x"898B8C8D", x"8C8C8D8D", x"91908F90", x"91918F8E", x"8F8F8F8E", x"8D8C8C8D", x"88868585", x"84807C79",
									 -- x"7A7D8285", x"837F7D7F", x"8281807D", x"7B7A7A7B", x"7E7C7B7C", x"7E7E7C7A", x"7F818483", x"807B7978",
									 -- x"78777A7C", x"7B7E7E79", x"7B7E7C7D", x"7B787C7A", x"7A7F7F7E", x"81828185", x"83848484", x"83838689",
									 -- x"8C868485", x"85878884", x"86898984", x"84888986", x"8B89888A", x"8D8E8D8B", x"8B8A8F8F", x"8E8E8989",
									 -- x"8D8C8B8D", x"8E8E8E8E", x"908F8D8C", x"8C8C8C8B", x"8C8C8A8A", x"8C8A898D", x"8A888A8B", x"8B8D8D88",
									 -- x"8B8A888C", x"8A888C88", x"8D8A8A8C", x"8A848589", x"86838387", x"86828285", x"88858184", x"8A8A8A8E",
									 -- x"8A8B8A8C", x"90909093", x"9193908E", x"91929091", x"9595989C", x"9C9B9DA2", x"AAA6A5AB", x"B0AAA6AC",
									 -- x"A4A7AEAB", x"A7A7A5A7", x"A6ABADAC", x"ACACAFB5", x"ADB1B3B0", x"AEAFAFAE", x"B1B0B0B1", x"B2B2B1B0",
									 -- x"ADABABAE", x"AFACABAC", x"B1B3B1B0", x"B4B5B4B3", x"B5B4B5B7", x"B6B2B1B3", x"B4B2AFAD", x"ACACAFB3",
									 -- x"B1B2B3B4", x"B5B6B6B6", x"B6B4B5B6", x"B1B0B3B4", x"B4B3B3B4", x"B5B5B7B9", x"BBB9B7B7", x"B8B9B9B9",
									 -- x"BEBBBCBD", x"BBBDC0BF", x"C0BFBEBD", x"BCBCBBBA", x"BCBBBABA", x"BCBDBCBC", x"BDBCBAB9", x"BABBB9B5",
									 -- x"9AA09F9C", x"9E9F9F9F", x"A3A3A4A5", x"A6A8AAAB", x"ADAEAFB0", x"AFADAEAF", x"B2B1AFAE", x"AEAFB0B1",
									 -- x"AFB0B1B2", x"B2B2B3B4", x"B5B5B5B6", x"B7B8B9BA", x"BDBDBDBF", x"C2C3C3C2", x"C2C2C4C5", x"C6C6C6C5",
									 -- x"C8C7C6C7", x"C8C8C6C5", x"C4C6C6C5", x"C6C7C7C5", x"C5C4C2C1", x"C2C3C5C6", x"C3C1C0BF", x"C0C1C2C3",
									 -- x"C1C1C1C1", x"C0C0C0BF", x"BFC1C1C0", x"C0C1C2C2", x"BFC3C4C3", x"C3C6C7C5", x"C8C8C8C8", x"C7C7C7C7",
									 -- x"C9C8C8C9", x"CCCFD0D0", x"CFD0D0CF", x"CECDCCCC", x"CBCAC8C7", x"C6C6C6C5", x"C6C5C4C5", x"C4C3C3C4",
									 -- x"C3C3C4C3", x"C2C1C0BF", x"C1C0BFC0", x"C1C1C2C2", x"C1C1C2C2", x"C3C3C4C5", x"C2C3C3C4", x"C5C5C5C5",
									 -- x"C6C8C9C8", x"C8CACAC8", x"C7C7C6C7", x"C7C6C7C7", x"CACAC9C7", x"C7C7C5C3", x"C4C3C4C4", x"C4C3C3C3",
									 -- x"C5C4C3C2", x"C0C0C0C0", x"C0C0C0C0", x"C0BFBEBD", x"BFBFBFBE", x"BCBCBCBD", x"BFC0C0BF", x"BDBCBBBB",
									 -- x"BBBAB9B8", x"B6B3B2B4", x"B3B1ADA9", x"A6A3A09F", x"98969596", x"97989898", x"95969490", x"8E8E8E8D",
									 -- x"8B8C8D8D", x"8D8D8D8D", x"93929191", x"92919190", x"90909090", x"8F8E8E8E", x"8B868383", x"817E7E80",
									 -- x"7D818688", x"857F7C7D", x"8281807E", x"7D7B7B7B", x"7F7D7C7D", x"7F808080", x"7F838687", x"84807E7E",
									 -- x"7E7D7F80", x"7E7F7F7A", x"7E807B7D", x"7D7B807E", x"7D808283", x"85858483", x"83858685", x"82818488",
									 -- x"8B868282", x"84878784", x"84888986", x"85888988", x"8B89888A", x"8C8B8A8A", x"89888B8E", x"8E8A8789",
									 -- x"8B8B8C8D", x"8E8F9091", x"91908D8C", x"8D8F908F", x"8E8F8E8E", x"8F8D8B8F", x"898A8B8A", x"8B8D8C86",
									 -- x"8B89878C", x"8A868B89", x"8C898888", x"86828387", x"89858383", x"84838689", x"8C898483", x"898B8A8D",
									 -- x"8A8D8D91", x"96918D93", x"8C908E8B", x"8E91908F", x"9494969A", x"9C9C9EA1", x"A3A3A4AA", x"AEAAA8AC",
									 -- x"A7ABAFAD", x"A9A8A7AA", x"A8AAA6A6", x"AEB0ADB0", x"AEB2B3B1", x"AEAEAFAF", x"B0AFAEAF", x"B0B1B0AE",
									 -- x"ADACADAE", x"AFAEADAD", x"B0B3AFAE", x"B3B3B0B3", x"B4B4B4B5", x"B5B3B2B2", x"B2B0ADAB", x"AAABAEB1",
									 -- x"B1B2B3B5", x"B6B6B6B6", x"B3B1B4B4", x"B0B0B3B2", x"B3B2B2B2", x"B3B4B5B7", x"B6B6B6B6", x"B7B8B8B8",
									 -- x"BEBCBDBE", x"BBBCBFBE", x"C3C0BEBC", x"BCBDBDBE", x"BCBAB9BA", x"BBBCBBB9", x"BBBCBAB8", x"B8BBBBB7",
									 -- x"969D9E9C", x"9E9F9E9F", x"A2A3A3A4", x"A4A7AAAC", x"AAACAEAE", x"ADADAEAE", x"ACACADAF", x"B0B1B3B3",
									 -- x"B3B2B0B0", x"B1B2B3B4", x"B3B4B6B7", x"B9B9BABA", x"BCBCBDBF", x"C2C3C3C2", x"C3C4C5C6", x"C6C6C6C6",
									 -- x"C9C8C8C9", x"CAC9C7C4", x"C5C6C6C5", x"C5C6C6C5", x"C4C4C3C2", x"C2C2C3C3", x"C2C1C0C0", x"C1C1C1C0",
									 -- x"C0C0C0C0", x"C0C0C0C0", x"BEC0C0BE", x"BEC0C1C1", x"BFC2C4C1", x"C1C5C5C3", x"C5C5C6C6", x"C6C6C6C5",
									 -- x"C8C7C7C9", x"CCCFD0D0", x"CFD0D0D0", x"CECDCDCD", x"CAC9C7C7", x"C7C6C6C6", x"C4C3C3C5", x"C5C3C2C3",
									 -- x"C3C3C2C2", x"C1C1C0C0", x"C1C0C0C0", x"C0C1C1C1", x"BFBFC0C0", x"C0C1C2C3", x"C1C2C3C3", x"C4C4C5C5",
									 -- x"C6C7C7C6", x"C6C7C8C7", x"C4C5C5C5", x"C5C5C5C4", x"C4C7C9C7", x"C5C5C4C2", x"C3C3C3C3", x"C3C3C2C2",
									 -- x"C3C2C1C0", x"C0C0C0C0", x"C1C0BFBF", x"BEBEBEBE", x"BDBEBDBC", x"BBBABABB", x"BDBDBEBF", x"BDBBBAB9",
									 -- x"BAB8B7B6", x"B4B2B1B2", x"B1AEAAA7", x"A4A3A2A1", x"9B9A9897", x"97989998", x"95959290", x"9191908D",
									 -- x"8C8D8E8E", x"8D8D8E8E", x"90909192", x"94959696", x"8F909090", x"8F8E8D8D", x"8E898584", x"817F8085",
									 -- x"82858889", x"86817F80", x"80808080", x"807E7D7C", x"7F7F7F7F", x"7F808386", x"81848788", x"87858585",
									 -- x"81818384", x"8183837E", x"81837E80", x"807E817F", x"81818385", x"8483817F", x"80838685", x"82818386",
									 -- x"8483807F", x"83848484", x"84888A88", x"86888887", x"8A898889", x"88868688", x"8888898D", x"8C878789",
									 -- x"878A8D8D", x"8D8E9294", x"91918E8C", x"8D919290", x"8E8F8D8C", x"8E8B8A8E", x"8E908F8B", x"8B8B8783",
									 -- x"87858389", x"86838887", x"8A8A8987", x"84848586", x"86868481", x"81858787", x"888A8581", x"868B8B8A",
									 -- x"8A8D8C8F", x"928D8A90", x"898E8C89", x"8D908E8E", x"9695969B", x"9EA09F9F", x"9EA5A7A8", x"AAAAA9AB",
									 -- x"ABACACAC", x"AAA8A9AA", x"ACADA7A6", x"ACACA8AA", x"B1B4B5B3", x"B0B0B1B1", x"AFAFB0B0", x"AFAFAFAE",
									 -- x"ACAFAFAC", x"ADB0AFAB", x"AFB1ADAB", x"B0AFADB2", x"B0B1B2B2", x"B2B2B1B0", x"AFAEADAC", x"ABACAEAF",
									 -- x"B1B2B3B4", x"B5B5B5B5", x"B0B2B4B2", x"AFB2B4B0", x"B2B2B2B2", x"B2B4B5B5", x"B4B6B8B9", x"B8B7B8B9",
									 -- x"BBBABDBE", x"BBBBBDBB", x"C2C0BEBD", x"BCBCBCBC", x"B8B8B7B8", x"B9BAB9B8", x"BABBBAB7", x"B8BBBAB6",
									 -- x"939A9C9D", x"A0A09FA1", x"A1A2A3A3", x"A4A6A9AC", x"A9ABADAD", x"ADAEAFAE", x"ABADB0B3", x"B4B3B2B1",
									 -- x"B6B3B0B1", x"B1B2B3B4", x"B3B5B7B9", x"BABBBBBA", x"BCBCBEC0", x"C3C5C4C3", x"C4C5C5C6", x"C6C7C7C7",
									 -- x"C8C9CACB", x"CBCAC7C5", x"C6C7C7C6", x"C5C7C6C5", x"C4C4C5C5", x"C4C2C0BE", x"C1C1C1C2", x"C2C2C0BF",
									 -- x"BEBEBEBF", x"BFC0C1C1", x"BEC0BFBC", x"BCBFC0C0", x"BEC1C1C0", x"C0C3C4C3", x"C3C3C3C4", x"C5C5C4C4",
									 -- x"C6C6C7C9", x"CBCECFCF", x"CECFD0CF", x"CECDCCCC", x"CAC7C6C7", x"C7C6C6C7", x"C3C2C2C5", x"C5C4C2C2",
									 -- x"C5C3C0BF", x"BFBFC1C3", x"C1C1C1C0", x"C0C2C2C0", x"BFC0C0C0", x"C0C0C1C2", x"C0C1C2C2", x"C3C3C4C4",
									 -- x"C5C4C4C4", x"C5C5C5C4", x"C2C3C3C3", x"C3C4C4C3", x"C2C6C8C7", x"C5C4C3C2", x"C3C4C3C2", x"C1C2C3C2",
									 -- x"C1C1C0C0", x"C0C0C0C0", x"C1C0BFBE", x"BDBDBDBE", x"BABBBBBA", x"B9B9BABA", x"BABABCBD", x"BCB9B8B8",
									 -- x"BAB8B6B6", x"B4B2B1B2", x"AEACA9A6", x"A4A3A2A1", x"9F9F9D9A", x"98989898", x"96959392", x"9394928F",
									 -- x"8E8F8F8F", x"8E8E8F8F", x"91929394", x"95959595", x"8D8E908F", x"8E8C8B8B", x"8D8B8987", x"84818284",
									 -- x"8787898A", x"89868587", x"82828383", x"8382807F", x"80818281", x"80808487", x"82838586", x"86868686",
									 -- x"7F7F8283", x"81838581", x"83868385", x"8480827E", x"87838586", x"8280817E", x"80828484", x"83828384",
									 -- x"81848281", x"86858486", x"83878988", x"86868584", x"88888886", x"85848586", x"898A888C", x"8A848787",
									 -- x"888D8F8D", x"8A898C8E", x"90908D8B", x"8C8F8F8B", x"8B8B8887", x"8987868A", x"8B8E8B87", x"89878484",
									 -- x"86858488", x"85838A88", x"86888885", x"84848484", x"80838380", x"7F82817D", x"7F85827E", x"83898987",
									 -- x"8A8C8B8B", x"8B898A90", x"8D908E8D", x"90918F90", x"97969699", x"9C9D9D9C", x"9EA7A9A6", x"A6A7A7A8",
									 -- x"AAABA7A9", x"A9A5A8A7", x"A8ACABA9", x"A9A9AAAE", x"B1B2B2B1", x"B0B0B0B0", x"ADAEAFAE", x"ADACACAC",
									 -- x"AAAEADA8", x"A9AEAEA9", x"ADADABAB", x"ADADADB0", x"B0B2B2B1", x"B1B3B3B0", x"ADAEAEAD", x"AEAFAFAE",
									 -- x"B1B2B2B2", x"B2B3B3B3", x"B1B3B5B2", x"AEB2B4AF", x"B3B3B3B2", x"B2B4B5B5", x"B3B6B9B9", x"B7B6B7B8",
									 -- x"BCBBBEBF", x"BDBDBEBB", x"BEBEBEBE", x"BDBBB8B6", x"B4B5B6B7", x"B8B8B9B9", x"B9BABAB9", x"B9B9B8B5",
									 -- x"95989A9D", x"A1A09FA3", x"A0A1A2A3", x"A3A4A8AA", x"AAACADAD", x"AEB0B0AE", x"AFB1B2B4", x"B4B2B1AF",
									 -- x"B3B2B2B3", x"B2B2B3B6", x"B5B6B8B9", x"BABBBBBB", x"BCBDBEC1", x"C5C6C6C5", x"C5C5C5C6", x"C7C8C9CA",
									 -- x"C8C9CBCC", x"CBC9C8C8", x"C6C7C7C5", x"C5C6C6C5", x"C3C4C4C3", x"C2C1C0BF", x"C0C0C1C2", x"C2C1C0BF",
									 -- x"BEBEBEBE", x"BEBFBFC0", x"BDBFBEBA", x"B9BDC0BF", x"BEBEBEBE", x"BEC0C2C3", x"C3C2C3C4", x"C5C5C3C2",
									 -- x"C4C5C8CA", x"CBCCCDCE", x"CDCECECE", x"CDCCCBCB", x"C9C7C5C6", x"C7C5C5C6", x"C5C3C2C4", x"C5C3C2C3",
									 -- x"C3C1C0C0", x"C0BFBFC1", x"BFC0BFBE", x"BFC2C2C0", x"C1C2C2C2", x"C1C1C2C3", x"C0C1C1C2", x"C2C2C2C2",
									 -- x"C3C2C2C2", x"C3C3C2C1", x"C0C1C2C1", x"C1C3C3C2", x"C2C4C5C4", x"C3C4C3C1", x"C2C3C2BF", x"BFC1C2C2",
									 -- x"C1C1C1C1", x"C1C1C1C0", x"C0BFBFBE", x"BDBCBCBC", x"B9BABAB9", x"B9B9B9BA", x"B9B8B8BA", x"B9B7B7B9",
									 -- x"B8B6B4B4", x"B3B2B1B3", x"ADACA9A7", x"A5A3A1A0", x"A1A19F9B", x"99999998", x"97979593", x"93959593",
									 -- x"90919191", x"90909091", x"96969796", x"95939291", x"8D8E8F8F", x"8E8C8A89", x"898B8B87", x"84838485",
									 -- x"8A898A8B", x"8C8B8B8C", x"89888786", x"86858483", x"82848586", x"85858687", x"84848586", x"88888786",
									 -- x"86868889", x"87898C89", x"8B8E8A8C", x"8A878A89", x"89838687", x"82818584", x"84838383", x"84838282",
									 -- x"82858384", x"89878284", x"81858887", x"85858686", x"87888783", x"84878886", x"878B878A", x"87828785",
									 -- x"878B8C8A", x"87868787", x"8C8D8B89", x"8A8D8B86", x"89898687", x"8A888688", x"86888482", x"87858288",
									 -- x"87888788", x"84848A86", x"81818385", x"837F7E80", x"7D7E807F", x"7E7D7A78", x"7D828281", x"84868586",
									 -- x"86888B8A", x"87898D8E", x"8D8E8D8E", x"92918F92", x"95969797", x"97999C9E", x"9EA4A4A3", x"A4A4A4A7",
									 -- x"A6A8A3A8", x"A7A2A6A5", x"A5A6AAAB", x"A8AAAFB1", x"AFAEADAD", x"AEAEAEAD", x"ABABACAB", x"AAA9A9A9",
									 -- x"AAAAA8A6", x"A6A9A9A8", x"AAA8AAAC", x"ABAAACAC", x"B0B2B2B0", x"B0B3B2AE", x"ACADADAC", x"ACAFAFAD",
									 -- x"B0B0AFAF", x"AFB0B0B1", x"B3B1B3B2", x"AFB0B1AF", x"B1B2B1B0", x"B1B4B5B5", x"B2B4B5B5", x"B5B5B6B7",
									 -- x"BFBCBEC0", x"BFC0C0BC", x"BDBDBDBD", x"BCBAB8B6", x"B4B6B8B8", x"B7B6B7B8", x"B8B8B9BB", x"BBB9B6B6",
									 -- x"9696969A", x"9E9C9BA0", x"9FA1A2A2", x"A2A3A6A8", x"ACADAEAD", x"AFB2B1AE", x"AFAFAEAE", x"AFB0B1B2",
									 -- x"AFB0B2B4", x"B3B2B4B9", x"B7B8B8B9", x"BABABBBB", x"BBBCBEC1", x"C5C7C6C5", x"C5C5C5C6", x"C7C9CACC",
									 -- x"C8C9CBCB", x"CAC9C9C9", x"C5C6C5C4", x"C4C5C6C5", x"C3C2C0BE", x"BEBFC1C2", x"BFBFBFC0", x"C0C0BFBE",
									 -- x"C0BFBEBD", x"BDBDBDBD", x"BDBFBDB8", x"B8BCBFBF", x"BDBCBCBD", x"BDBEC0C3", x"C3C3C3C4", x"C4C4C2C1",
									 -- x"C2C5C8CA", x"CBCBCCCD", x"CBCCCDCD", x"CCCBCACA", x"C9C6C5C6", x"C6C5C5C6", x"C8C5C3C3", x"C4C3C3C4",
									 -- x"BFBFC1C4", x"C3C0BDBE", x"BCBEBEBC", x"BEC1C1BF", x"C1C1C1C1", x"C0C0C1C2", x"C1C1C1C1", x"C1C1C1C0",
									 -- x"C2C1C0C1", x"C2C2C0C0", x"BFC1C1C0", x"C0C3C3C1", x"C3C3C2C1", x"C2C3C1BF", x"C0C1C0BD", x"BDC0C2C1",
									 -- x"C1C2C2C2", x"C2C2C1C0", x"BFBFBFBE", x"BDBCBBBA", x"BABBBAB9", x"B8B8B8B9", x"B8B7B6B7", x"B7B6B7BA",
									 -- x"B6B4B2B2", x"B2B1B1B2", x"ADACABA9", x"A7A4A09E", x"9FA09E9A", x"99999A98", x"96969591", x"90929494",
									 -- x"92929292", x"91919292", x"96979797", x"95939191", x"8E8F9090", x"8F8C8A89", x"868A8A85", x"82858888",
									 -- x"8C8A8A8C", x"8D8D8C8C", x"8F8D8A88", x"88878685", x"84858789", x"8A8A8988", x"8988898B", x"8E8E8D8B",
									 -- x"8C8B8D8C", x"898B8D8A", x"8C8D8887", x"86868D8E", x"86808486", x"81828989", x"89868483", x"8383817F",
									 -- x"80848282", x"89867E7E", x"80848686", x"8586898B", x"86878581", x"848A8B87", x"848A8587", x"84808784",
									 -- x"7F838585", x"86888988", x"88898987", x"8A8D8A84", x"8B8B888A", x"8E8D898B", x"88888382", x"87838189",
									 -- x"878A8785", x"81818680", x"817D8086", x"847C7A7F", x"7E7C7C7F", x"7E7A787A", x"81848586", x"87838185",
									 -- x"7F838A8B", x"86898E89", x"8887878A", x"8F8D8C91", x"96989A98", x"97999FA4", x"9C9D9C9F", x"A3A2A2A8",
									 -- x"A2A6A2A8", x"A69FA5A3", x"A9A4A7AA", x"A8ACB0AC", x"B0ADACAD", x"AFAFAEAD", x"ABAAAAAA", x"AAA9A8A7",
									 -- x"ABA8A5A6", x"A6A5A6A8", x"A7A3A8AD", x"A9A8AAA8", x"ADB0AFAC", x"ADB0AFAA", x"ACADABA9", x"AAADAEAC",
									 -- x"AFAEADAD", x"ADAEAFB0", x"B4AEAFB2", x"AFADAEB0", x"AEAFAFAE", x"AFB2B4B3", x"B3B2B2B3", x"B5B8B9B9",
									 -- x"BEBABBBC", x"BCBEBFBB", x"BFBDBBBA", x"BABABABA", x"B7B9BBBA", x"B7B5B5B7", x"B7B6B8BD", x"BDB9B7B8",
									 -- x"94969A9D", x"9C9A9CA0", x"9F9E9FA0", x"A2A4A3A3", x"A8ABADAD", x"ADB0B1B0", x"ACB0B3B3", x"B0AEB0B2",
									 -- x"B1B1B4B6", x"B4B2B3B7", x"B9B9B8B8", x"B8BABDBF", x"C1C0C0C2", x"C4C5C5C5", x"C5C6C7C9", x"CACAC9C9",
									 -- x"CBC9C8C7", x"C8C9C9C9", x"C6C5C4C4", x"C5C4C3C1", x"C2C4C3BF", x"BDBEC0C0", x"C3C1C0C1", x"C2C1BEBB",
									 -- x"BBBCBDBE", x"BEBDBCBB", x"B7B8B9BA", x"BABABABA", x"BABABCBE", x"C0C1C0BF", x"C0C1C2C2", x"C1C0C1C2",
									 -- x"C5C7C8C8", x"C9CCCECE", x"CAC9C8C8", x"C9C8C7C6", x"C5C6C6C6", x"C5C5C6C6", x"C6C5C4C3", x"C2C1BFBD",
									 -- x"C2C1C0C0", x"BFBEBDBD", x"BDBEBEBD", x"BEC1C0BE", x"BEC0C1C0", x"C0C0BFBE", x"BDBFC0C1", x"C0C0C1C1",
									 -- x"C0C0C0BF", x"BFBFBFBE", x"C1C0BFBE", x"BEBEBFBF", x"BEBEBFBF", x"BFBFBFBE", x"BFBEBEBF", x"C0BFC0C1",
									 -- x"BFBFBFC0", x"C0C1C2C2", x"BFBFBEBD", x"BCBBBABA", x"B8BABCBB", x"B8B6B6B8", x"B8B8B7B6", x"B5B4B4B3",
									 -- x"B6B4B2B2", x"B2B2B0AE", x"ACA9A7A5", x"A5A4A19E", x"A09E9C99", x"9898999B", x"98979594", x"93939394",
									 -- x"91919191", x"92939597", x"99959497", x"97928E8D", x"92908E8E", x"8E8E8C8A", x"858A8B89", x"8C8C8A8B",
									 -- x"8C8C8B8D", x"9193928F", x"8B8D8D8C", x"8A888888", x"888B8D8B", x"898A8C8C", x"8D8E8E8D", x"8E90918F",
									 -- x"9192908F", x"8E8F8E8C", x"90908E8A", x"8A8D9091", x"8A878885", x"85888486", x"8A878587", x"87858281",
									 -- x"89888787", x"8785827F", x"7F848682", x"8084898B", x"88858382", x"83858686", x"85858C8C", x"83828684",
									 -- x"84848182", x"88868287", x"86888988", x"888A8A8A", x"898B8C8A", x"88888785", x"84838487", x"87838181",
									 -- x"82848582", x"81818180", x"827E7D80", x"83807C79", x"7A7A7F81", x"7C767575", x"80818384", x"83828386",
									 -- x"86858688", x"87858588", x"888A8B8B", x"898A8C8E", x"90969896", x"969A9E9E", x"A09E9D9E", x"9FA0A4A8",
									 -- x"A2A4A8A6", x"A1A3A8AA", x"A6A4A7AD", x"ACA8AAB1", x"A8A9A9A9", x"AAAAA9A9", x"A5A7A8A6", x"A6A7A8A6",
									 -- x"A8A19FA5", x"A7A4A3A7", x"A7A5A6AA", x"AAA7A6A8", x"ADABAAAC", x"ADACAAAA", x"A8A9AAAA", x"ABACACAB",
									 -- x"AAACACAB", x"ABADAEAC", x"ABAAABAD", x"AAA8ABB2", x"B2AFAFB1", x"B1B2B2AD", x"B0B4B5B3", x"B5BABBB9",
									 -- x"C1C0BDBA", x"BABDBEBD", x"BCBBBAB9", x"B9B9BABA", x"B8B9B7B4", x"B5B9B9B6", x"B9B9B8B8", x"BABCBCBA",
									 -- x"9696999B", x"9C9A9B9D", x"A09F9E9E", x"A0A2A4A4", x"A7A9ABAB", x"ACAFB0B0", x"B0B2B4B3", x"B1AFB0B1",
									 -- x"B5B4B5B6", x"B6B5B4B6", x"B7B8B8B9", x"BABCBEC0", x"C2C2C2C4", x"C5C5C4C4", x"C6C7C8C9", x"C9C9C9C9",
									 -- x"CAC9C8C7", x"C7C7C7C8", x"C7C6C6C6", x"C7C6C4C2", x"C3C4C3C0", x"BFC1C2C1", x"C1BFBEBE", x"BEBEBEBC",
									 -- x"BCBCBCBC", x"BCBBBAB9", x"B7B7B7B8", x"B9BABBBB", x"BCBBBBBA", x"BBBCBDBE", x"BFC0C1C1", x"C1C0C1C1",
									 -- x"C3C4C5C4", x"C4C6C8C8", x"C9C8C7C7", x"C7C7C7C6", x"C6C6C6C6", x"C5C4C5C5", x"C5C4C3C3", x"C2C1C0BF",
									 -- x"BFC0C0C0", x"BFBEBDBC", x"BCBDBDBC", x"BDC0BFBD", x"BCBEBEBD", x"BDBEBEBC", x"BDBEBFC0", x"C0C0C0C0",
									 -- x"BEBEBDBD", x"BCBDBDBD", x"BFBEBEBD", x"BDBDBEBE", x"BBBCBDBD", x"BEBDBDBC", x"BDBCBCBD", x"BDBCBDBF",
									 -- x"BEBEBFBF", x"C0C1C1C2", x"BFBEBCBA", x"B8B7B6B5", x"B6B9BBBA", x"B7B6B7B8", x"B7B7B6B6", x"B5B5B4B4",
									 -- x"B3B2B1B1", x"B2B1AFAD", x"ADAAA7A6", x"A5A4A2A0", x"9F9E9D9B", x"9A999999", x"97969594", x"94949596",
									 -- x"93939393", x"93949697", x"99969495", x"95939190", x"8E8E8E8F", x"908F8B89", x"868B8B8A", x"8D8E8C8E",
									 -- x"90909193", x"97989592", x"92929291", x"8F8D8E8F", x"8C8D8D8C", x"8C8D8D8C", x"9191908F", x"91939494",
									 -- x"95969594", x"94959593", x"93949494", x"92919090", x"918C8D89", x"898D8A8D", x"8A888787", x"87868687",
									 -- x"85848485", x"86868482", x"80858682", x"7F818484", x"85858484", x"84848483", x"87828485", x"8182837E",
									 -- x"85848284", x"88878688", x"8A8C8C8A", x"89898886", x"85868788", x"87878687", x"84848485", x"827F7E80",
									 -- x"807F7D7E", x"82868581", x"7E7C7C7F", x"807E7B7A", x"77777778", x"7775767A", x"767B8286", x"847F7D7F",
									 -- x"87848384", x"84828282", x"83858687", x"87898B8E", x"898E9395", x"9597999A", x"9F9FA0A0", x"A1A2A5A6",
									 -- x"A09EA0A3", x"A3A5A9A8", x"A8A6A7AB", x"A9A4A6AC", x"AAA9A9A9", x"A9A7A4A2", x"A1A4A5A3", x"A3A4A6A5",
									 -- x"A4A0A0A3", x"A3A0A0A3", x"A2A2A4A6", x"A6A6A8AA", x"ACAAA9AA", x"AAA8A8A9", x"A8A8A8A8", x"A8A7A4A2",
									 -- x"A7A9AAAA", x"AAADAEAE", x"B0ACABAE", x"AFADABAC", x"ABACB1B2", x"ADADB2B3", x"B0B2B4B4", x"B6B9BAB9",
									 -- x"BBBCBBB9", x"B7B8B7B5", x"B7B8B9B8", x"B7B7B9BA", x"B6B8B8B7", x"B6B7B9BA", x"B5B7B7B8", x"BABBBAB7",
									 -- x"97969799", x"9B9A9A9A", x"A09F9E9F", x"A1A3A4A5", x"A5A8A9AA", x"ABAEB0B0", x"B1B2B3B3", x"B2B1B1B1",
									 -- x"B5B4B3B5", x"B6B5B3B3", x"B5B7B8BA", x"BCBDBFC1", x"C1C3C5C6", x"C6C5C5C5", x"C7C8C8C9", x"C9C9C9C9",
									 -- x"C8C9C9C7", x"C6C5C6C7", x"C6C6C6C7", x"C8C7C5C2", x"C2C2C1BF", x"C0C1C0BF", x"BEBDBCBB", x"BBBCBDBE",
									 -- x"BFBFBEBD", x"BCBBBAB9", x"B7B7B6B6", x"B7B9BBBC", x"BABBBAB9", x"B8B9BBBD", x"BEBEBFC0", x"C1C1C1C0",
									 -- x"C2C4C4C3", x"C2C4C6C6", x"C8C7C6C5", x"C6C6C6C5", x"C6C6C6C6", x"C4C4C4C4", x"C4C3C2C1", x"C1C1C1C0",
									 -- x"BDBEBFBF", x"BFBDBCBB", x"BDBDBDBC", x"BDBFBFBE", x"BCBDBDBC", x"BCBDBDBC", x"BDBDBEBF", x"BEBEBFBF",
									 -- x"BDBDBCBC", x"BCBCBDBD", x"BDBDBDBD", x"BCBCBBBB", x"B8B9BABB", x"BBBBBABA", x"BABABBBC", x"BBBABBBE",
									 -- x"BCBCBDBE", x"BEBFBFC0", x"BEBCBAB8", x"B6B4B4B3", x"B4B7B9B9", x"B7B6B7B9", x"B8B7B6B5", x"B4B4B3B3",
									 -- x"B0AFB0B0", x"B1B0AEAB", x"ACAAA8A5", x"A3A2A2A2", x"9F9F9E9E", x"9C9B9998", x"98979695", x"95959697",
									 -- x"95959595", x"94959596", x"97979695", x"95969491", x"8D8D8E8F", x"90908D8B", x"8A8E8D8C", x"8F909092",
									 -- x"9394969A", x"9D9D9A97", x"96969593", x"91909193", x"92929090", x"9192918E", x"92929190", x"92969897",
									 -- x"9B9B9A98", x"97989694", x"93929395", x"938D8A8B", x"938E8D89", x"888C8A8D", x"8D8B8987", x"84838588",
									 -- x"83828284", x"85868584", x"83868581", x"7E808281", x"82848585", x"84828180", x"85807F7F", x"7E7F807C",
									 -- x"85818285", x"86878886", x"85868787", x"87888785", x"85848486", x"86838285", x"83838382", x"7E7C7D80",
									 -- x"827F7C7C", x"7F82807C", x"7B7B7C7C", x"7B787676", x"787A7573", x"7877777E", x"777A7D7E", x"7B797C81",
									 -- x"827F7D7E", x"81828281", x"81828385", x"878A8C8D", x"8A8C9195", x"9695979A", x"999D9F9E", x"9FA1A2A0",
									 -- x"A29EA0A4", x"A2A1A2A2", x"A09FA1A6", x"A7A5A8AD", x"ABAAA9A9", x"A8A6A29E", x"A0A2A3A2", x"A1A3A5A7",
									 -- x"A1A2A3A2", x"A0A09FA0", x"A0A2A3A2", x"A1A2A4A5", x"A9A8A8A8", x"A7A5A6A9", x"A6A6A7A8", x"A9A7A4A2",
									 -- x"A4A7A9A8", x"A8AAADAE", x"B0ACABAD", x"AEABAAAA", x"B0ACACAE", x"ADAEAFAC", x"AEAEAFB3", x"B5B5B6B8",
									 -- x"B7BABBBA", x"B8B6B5B4", x"B4B6B8B7", x"B5B4B6B8", x"B4B6B8B8", x"B6B4B7BC", x"B3B5B6B7", x"BABBB9B6",
									 -- x"94959698", x"9898999A", x"9D9EA0A3", x"A5A5A5A5", x"A6A7A9AA", x"ABADAFB0", x"B0B0B0B0", x"B1B2B2B1",
									 -- x"B4B3B4B4", x"B5B4B3B3", x"B5B7B8BA", x"BCBEC0C2", x"BFC2C5C5", x"C5C6C7C7", x"C8C8C8C9", x"C8C8C8C8",
									 -- x"C7C8C9C7", x"C5C5C6C8", x"C4C4C5C6", x"C7C6C4C2", x"C2C1BFBF", x"C0C0BFBD", x"BDBDBCBB", x"BABBBDBE",
									 -- x"BFBFBEBD", x"BCBBBAB9", x"B7B7B6B6", x"B7B8BABB", x"B7B9BBBB", x"B9B9BABC", x"BEBDBDBE", x"C0C2C1C0",
									 -- x"C1C3C5C4", x"C4C6C6C6", x"C7C6C5C4", x"C4C4C5C5", x"C5C6C6C5", x"C4C3C3C4", x"C4C2C1C0", x"C1C1C0C0",
									 -- x"BDBDBDBE", x"BDBDBCBC", x"BDBDBDBD", x"BDBEBFBF", x"BEBFBFBE", x"BDBEBEBC", x"BEBEBEBE", x"BDBDBDBD",
									 -- x"BDBCBCBC", x"BCBCBCBD", x"BCBCBCBC", x"BBBAB9B8", x"B8B8B8B8", x"B8B8B8B8", x"B9B9BBBC", x"BBB9BABD",
									 -- x"BABBBBBC", x"BDBDBEBE", x"BDBCB9B7", x"B5B5B5B5", x"B3B5B7B8", x"B7B7B9BA", x"B9B8B6B5", x"B3B2B1B1",
									 -- x"AEAEAFB0", x"B0AFACAA", x"AAA9A8A5", x"A3A1A1A1", x"9F9F9F9E", x"9E9C9A98", x"9B999896", x"95959696",
									 -- x"95959695", x"95959596", x"93979897", x"9797948E", x"908F8E8E", x"8F90908F", x"8E92908E", x"91939395",
									 -- x"9696989D", x"9F9E9C9A", x"98989795", x"93939495", x"97979594", x"95979593", x"93949393", x"95999A9A",
									 -- x"9D9E9D9B", x"9B9B9997", x"9D999799", x"96908E92", x"938E8E89", x"888B888B", x"8F8C8987", x"8585878A",
									 -- x"86858484", x"85858584", x"8586847F", x"7F838584", x"81838686", x"84828080", x"8080807F", x"7C7C7E7F",
									 -- x"837E8184", x"81838682", x"81828282", x"84878785", x"86838386", x"85808084", x"82828281", x"7F7E7F81",
									 -- x"81817F7C", x"7979797A", x"7A7C7C7B", x"78757577", x"7B7F7875", x"7C7A757B", x"7B7A7876", x"74757C84",
									 -- x"7D7B7B7D", x"80828181", x"80808183", x"86898B8B", x"908E8F93", x"93909398", x"959B9D9B", x"9B9F9F9B",
									 -- x"A0A0A5A7", x"9F9A9DA1", x"A4A3A5A7", x"A7A4A4A6", x"A9A8A7A7", x"A8A7A4A1", x"9EA0A1A0", x"9FA0A3A6",
									 -- x"9FA3A3A0", x"9EA09F9B", x"9CA1A39F", x"9D9FA1A1", x"A2A3A5A6", x"A3A1A3A6", x"A5A5A7A9", x"A9A7A5A5",
									 -- x"A3A5A7A7", x"A5A6A9AC", x"AAAAA9A8", x"A6A4A9AF", x"B3ABA9AC", x"ADAEADA9", x"AEABADB3", x"B4B2B3B7",
									 -- x"B5B8BABA", x"B8B7B7B8", x"B6B7B8B6", x"B4B3B3B4", x"B3B4B6B7", x"B4B1B3B8", x"B4B5B6B6", x"B8BABAB8",
									 -- x"92959796", x"95959799", x"9B9D9FA2", x"A4A5A5A5", x"A7A8A9AA", x"ABACAEB0", x"B0B0AFB0", x"B1B2B2B1",
									 -- x"B2B4B6B6", x"B5B4B5B6", x"B7B7B9BA", x"BBBEC0C2", x"BFC3C5C4", x"C3C5C7C7", x"C8C8C8C8", x"C8C8C7C7",
									 -- x"C5C7C8C8", x"C6C6C7C9", x"C5C4C4C4", x"C5C5C4C3", x"C4C2C1C1", x"C1C0BEBD", x"BDBEBEBD", x"BCBCBDBE",
									 -- x"BBBBBCBB", x"BAB9B7B6", x"B7B7B7B8", x"B8B8B9B9", x"B7B9BABA", x"B9B8BABB", x"BDBCBCBE", x"C0C1C1C0",
									 -- x"BFC2C4C4", x"C4C5C4C3", x"C5C5C4C3", x"C3C3C4C5", x"C4C5C5C4", x"C4C3C3C4", x"C4C3C1C0", x"C0C0BFBF",
									 -- x"BEBDBDBC", x"BCBCBDBD", x"BCBCBCBC", x"BCBCBDBF", x"BFC0C0BF", x"BEBEBEBC", x"BFBFBFBE", x"BCBBBBBB",
									 -- x"BBBAB9BB", x"BBB9B9BB", x"BABABBBB", x"BAB9B8B7", x"B9B8B7B6", x"B5B6B7B7", x"B8B8BABB", x"BAB9BABC",
									 -- x"BBBBBCBC", x"BDBDBDBD", x"BCBBB9B7", x"B5B4B4B4", x"B3B4B7B8", x"B8B8B9BA", x"BAB9B7B4", x"B1AFAEAE",
									 -- x"ADAEAEAF", x"AEADAAA9", x"A8A9A8A7", x"A4A2A0A0", x"9F9E9E9E", x"9D9C9A99", x"9B9A9896", x"95959696",
									 -- x"95959696", x"96969697", x"94979997", x"9797938E", x"91908F8E", x"8F8F9090", x"90949391", x"9496979A",
									 -- x"9B9A9B9F", x"A19F9D9D", x"9B9C9C9B", x"99989899", x"98999998", x"97989897", x"98999999", x"9A9C9C9A",
									 -- x"9C9E9F9F", x"A1A3A3A1", x"A29D9A9B", x"98939397", x"9491928E", x"8E908C8D", x"8D8A8788", x"8A8B8C8D",
									 -- x"89888786", x"86868585", x"84858481", x"81858684", x"81838585", x"83828181", x"7D7F807E", x"7E7C7D7F",
									 -- x"807D7F81", x"7D80827E", x"83848381", x"82848483", x"827F7F83", x"83808186", x"83828181", x"82828280",
									 -- x"7E7E7C7B", x"79797B7D", x"7B7C7D7B", x"7878797B", x"7B7F7774", x"7B797377", x"78767677", x"7676797C",
									 -- x"7B7D7F80", x"807F7E7D", x"7D7D7E80", x"83868889", x"8F8B8C8F", x"8E8B8D93", x"969B9D9A", x"9B9F9F9C",
									 -- x"9C9DA3A6", x"A19EA1A3", x"A4A5A7A9", x"AAA9A7A6", x"A7A5A4A4", x"A6A7A5A4", x"9C9D9E9E", x"9D9D9FA1",
									 -- x"9DA09F9A", x"9B9F9C95", x"969CA09E", x"9C9FA1A0", x"9C9FA2A3", x"A09D9DA0", x"A4A4A6A7", x"A4A0A1A4",
									 -- x"A1A3A5A4", x"A3A3A6A9", x"A7A7A7A6", x"A4A4A8AE", x"ABA9ACAE", x"ABAAAEB0", x"AFACAEB4", x"B6B4B4B9",
									 -- x"B4B5B6B6", x"B5B4B7B9", x"B9B8B6B6", x"B5B4B2B1", x"B4B2B2B5", x"B4B2B2B6", x"B6B6B4B3", x"B5B9BAB9",
									 -- x"91959795", x"93939597", x"9A9B9C9D", x"9EA1A4A6", x"A7A7A8A9", x"AAABADAF", x"B1B1B1B1", x"B2B2B1B0",
									 -- x"AFB3B5B5", x"B3B4B5B6", x"B7B8B9B9", x"BBBDC0C2", x"C1C4C4C2", x"C2C5C6C5", x"C7C7C8C8", x"C8C7C6C6",
									 -- x"C4C6C7C7", x"C6C6C7C9", x"C7C5C4C5", x"C5C6C4C3", x"C4C2C1C1", x"C0BEBDBC", x"BEBEBEBE", x"BEBDBDBD",
									 -- x"BABABABA", x"B9B8B7B6", x"B6B7B8B9", x"B9B8B8B7", x"BABAB9B8", x"B6B7B9BB", x"BCBCBDBE", x"C0C1C1C0",
									 -- x"C0C3C5C4", x"C4C4C3C1", x"C4C4C4C3", x"C2C2C3C4", x"C4C4C4C4", x"C3C3C3C3", x"C4C3C1C0", x"C0BFBEBD",
									 -- x"BEBDBCBB", x"BBBBBCBD", x"BAB9B9B9", x"B9B9BABD", x"BDBEBFBE", x"BDBDBCBA", x"BEBEBEBC", x"BBB9B9BA",
									 -- x"BCB9B9BB", x"BBB8B8BB", x"B7B7B8B9", x"B9B9B8B8", x"B7B6B5B4", x"B3B4B5B6", x"B7B6B7B9", x"B9B8B8B9",
									 -- x"BCBCBDBD", x"BDBDBCBC", x"BBBAB7B5", x"B3B2B1B1", x"B3B4B6B7", x"B8B9B9BA", x"BAB8B5B2", x"B0AEADAC",
									 -- x"ADADADAD", x"ACABA9A9", x"A9A9A8A8", x"A6A3A19F", x"9E9D9C9C", x"9D9D9B99", x"9A999796", x"95969697",
									 -- x"96969797", x"97979899", x"98999997", x"95959492", x"8F909191", x"91908F8E", x"92959493", x"979A9B9F",
									 -- x"A19FA0A3", x"A4A19FA0", x"9F9FA09E", x"9C9B9C9D", x"9A9B9B9A", x"999A9A99", x"9D9E9E9D", x"9D9D9C99",
									 -- x"9FA1A2A3", x"A4A6A6A4", x"9D9B9A9A", x"97939295", x"918F928F", x"90928D8F", x"8D898688", x"8A8A8989",
									 -- x"88888887", x"87878787", x"81848684", x"83858480", x"82828383", x"82828181", x"7E7E7B7B", x"807F7B7B",
									 -- x"7E7D7E7E", x"7C7E7F7C", x"8082817F", x"7E808181", x"827F7F80", x"7F7E7F82", x"85848281", x"8283817D",
									 -- x"807B7879", x"7D7E7D7C", x"7C7D7C79", x"77767675", x"797B7571", x"76777578", x"75737374", x"75747475",
									 -- x"767A7F80", x"807F7E7C", x"7B7C7D7F", x"82858789", x"8D8A8C90", x"908D8E92", x"969A9A99", x"999D9E9D",
									 -- x"9E9B9EA2", x"A3A4A49F", x"9B9EA1A5", x"A9ABAAA8", x"A4A3A2A1", x"A2A2A2A2", x"9C9B9C9E", x"9D9C9C9D",
									 -- x"9C9D9B97", x"989D9B95", x"979A9D9D", x"9C9D9D9D", x"9D9FA2A3", x"A09C9B9C", x"A0A0A2A4", x"A29FA0A4",
									 -- x"A0A0A1A2", x"A1A1A3A7", x"A7A6A5A6", x"A8A9A8A7", x"ACA7A8AC", x"ABABADAC", x"ADABADB3", x"B5B3B3B7",
									 -- x"B5B4B3B3", x"B2B2B4B8", x"B9B6B4B4", x"B5B5B3B1", x"B3B1B0B2", x"B4B5B5B5", x"B6B5B2B1", x"B3B7B8B8",
									 -- x"8F929493", x"92949696", x"9A9A9B9B", x"9C9EA1A4", x"A5A4A5A7", x"A8A9ABAE", x"B0B0B1B2", x"B2B1B0B0",
									 -- x"AEB1B3B2", x"B2B4B4B4", x"B6B7B8BA", x"BBBDBFC1", x"C1C4C4C2", x"C4C7C6C3", x"C5C6C7C8", x"C8C7C6C5",
									 -- x"C5C5C5C6", x"C6C6C7C7", x"C7C6C5C6", x"C7C6C4C2", x"C2C1C0C0", x"BFBCBBBD", x"BFBEBDBD", x"BEBEBDBC",
									 -- x"BCBAB9B7", x"B7B7B7B7", x"B5B6B7B8", x"B8B8B7B7", x"BBBAB9B8", x"B8B9BABB", x"BCBDBEBF", x"BFC0C0C1",
									 -- x"C1C3C4C4", x"C3C4C4C3", x"C3C4C4C4", x"C3C2C3C4", x"C4C4C4C4", x"C3C2C2C2", x"C3C2C1C0", x"C0BFBDBC",
									 -- x"BDBCBBBA", x"BABABBBB", x"B8B7B7B8", x"B7B7B9BC", x"B9BBBDBD", x"BDBDBBB9", x"BCBCBCBA", x"B9B8B8B9",
									 -- x"BDB9B9BB", x"BAB7B7BA", x"B6B6B7B7", x"B7B7B6B6", x"B2B2B2B2", x"B2B2B3B3", x"B6B5B5B7", x"B9B8B7B6",
									 -- x"BBBBBCBC", x"BCBBBAB9", x"B8B7B5B3", x"B2B0AFAF", x"B3B4B5B7", x"B7B8B8B8", x"B7B5B3B1", x"AFAEADAD",
									 -- x"ACABABAA", x"A9A9A9A9", x"A9A8A6A5", x"A5A3A09E", x"9C9B9B9C", x"9D9D9B99", x"99989795", x"95959696",
									 -- x"97979796", x"9697989A", x"9B9A9999", x"97959596", x"91929393", x"93929191", x"94989795", x"999B9DA0",
									 -- x"A4A2A3A7", x"A8A5A4A6", x"A2A2A2A0", x"9E9E9FA0", x"9F9F9E9C", x"9D9E9D9A", x"9FA09F9E", x"9E9F9E9C",
									 -- x"A2A4A4A4", x"A5A6A5A3", x"A1A09F9D", x"9A999999", x"908D908E", x"8E908C8D", x"8F8C8A89", x"88868484",
									 -- x"87878787", x"87868787", x"82868784", x"83848381", x"82828282", x"8281807F", x"7D807C7A", x"7F7D787A",
									 -- x"7A7D7C7A", x"7B7C7B7C", x"7A7D807E", x"7C7D7E7F", x"8382817F", x"7D7D7E7F", x"8484827F", x"7F807E7B",
									 -- x"827C7879", x"7B7A7877", x"7B7B7A78", x"7877736E", x"77777471", x"72747576", x"74727170", x"706F7174",
									 -- x"72767B7D", x"7F807D79", x"7C7D7F80", x"81838587", x"8A88898C", x"8D8D8F92", x"94959697", x"98999B9C",
									 -- x"9E9C9D9F", x"A1A5A39A", x"9E9F9F9F", x"A2A3A19D", x"A1A2A2A0", x"9E9D9D9E", x"9A999A9D", x"9E9C9A99",
									 -- x"9A9B9995", x"969A9A97", x"9A9A9B9C", x"9B9A9A9B", x"9D9EA1A2", x"A09C9B9C", x"9C9A9CA1", x"A2A09FA2",
									 -- x"A1A09FA0", x"A09FA0A3", x"A4A4A3A5", x"A7A8A7A5", x"AEA4A2A8", x"ACACAAA5", x"A9A9ABAF", x"B1B1B1B3",
									 -- x"B5B3B2B3", x"B3B1B2B4", x"B6B5B3B2", x"B3B3B3B2", x"B1B1B0B0", x"B2B5B5B4", x"B5B4B3B3", x"B4B7B7B5",
									 -- x"8D8F9090", x"93979897", x"989A9C9D", x"9D9E9FA1", x"A3A2A3A5", x"A7A7AAAD", x"ACAEB0B1", x"B1B0B0B0",
									 -- x"B0B2B2B2", x"B4B6B6B3", x"B4B6B8BB", x"BCBEBFC0", x"BFC3C4C3", x"C5C9C8C3", x"C4C5C7C8", x"C8C7C5C4",
									 -- x"C5C4C4C5", x"C6C6C5C5", x"C6C5C6C6", x"C7C6C3C1", x"C3C1C1C2", x"BFBCBDC0", x"BFBDBBBC", x"BDBEBDBC",
									 -- x"BBB9B6B4", x"B3B3B5B6", x"B4B5B6B7", x"B7B8B7B7", x"B9B9BABC", x"BDBDBCBB", x"BBBDBFBF", x"BFBFC0C1",
									 -- x"BFC1C2C1", x"C1C3C4C4", x"C2C3C4C4", x"C3C2C3C3", x"C5C5C5C4", x"C2C1C1C1", x"C2C1C1C0", x"C0BFBDBC",
									 -- x"BBBBBBBB", x"BABAB9B9", x"B8B7B7B8", x"B7B6B8BC", x"B7BABCBC", x"BDBDBBB9", x"BABABAB9", x"B7B7B8B8",
									 -- x"BBB7B7B9", x"B8B4B4B7", x"B7B7B7B6", x"B5B4B3B2", x"AEAFB0B1", x"B1B2B1B1", x"B7B5B4B7", x"BAB9B7B6",
									 -- x"B9B9B9BA", x"B9B8B7B6", x"B5B5B4B3", x"B2B1B0AF", x"B3B4B5B6", x"B7B7B7B7", x"B4B3B1AF", x"AEAEAEAF",
									 -- x"AAAAA9A8", x"A7A7A9AA", x"A8A6A3A2", x"A2A19F9D", x"9A9A9A9C", x"9D9D9A98", x"9A999795", x"94949494",
									 -- x"96969695", x"95959798", x"9A999A9D", x"9B969596", x"95959493", x"93949597", x"979B9997", x"999B9B9E",
									 -- x"A2A1A4A9", x"ABA9A8AB", x"A6A5A4A2", x"A0A0A2A4", x"A5A3A09F", x"A1A3A09C", x"A1A1A1A0", x"A1A3A3A2",
									 -- x"A2A4A5A6", x"A7A9A8A6", x"A3A3A09B", x"999B9C9D", x"94919390", x"90918D8E", x"918F8E8D", x"8A878789",
									 -- x"85868786", x"86858586", x"85888682", x"80838585", x"83828181", x"81817F7D", x"7B82817C", x"7C77767E",
									 -- x"767C7A77", x"7B7B787B", x"7A7F8281", x"7D7C7D7D", x"8182817E", x"7E808181", x"8283817E", x"7C7D7D7B",
									 -- x"7D7B7A79", x"77747477", x"76777879", x"7C7D7872", x"75757572", x"6F70716E", x"70717273", x"706D6E71",
									 -- x"7476797B", x"7D7E7973", x"7B7D7E7E", x"7D7E8183", x"85838181", x"83868B8E", x"93939497", x"9898999C",
									 -- x"999B9F9E", x"9DA3A39B", x"9C9D9D9C", x"A0A3A29F", x"A0A1A2A1", x"9E9C9B9C", x"9795979B", x"9D9B9795",
									 -- x"96989692", x"91959797", x"9996969A", x"9B9A9B9E", x"999A9C9E", x"9D9B9A9C", x"9D99999E", x"A19E9A99",
									 -- x"A3A09F9F", x"9E9D9DA0", x"9FA1A3A2", x"A0A1A5A9", x"A5A0A3A9", x"A8A7A9AA", x"A8A9ABAF", x"B1B1B2B2",
									 -- x"B1AFAFB2", x"B2B1B0B1", x"B5B4B3B2", x"B1B0B1B2", x"B0B2B1AE", x"AFB2B3B1", x"B4B5B6B6", x"B7B8B6B3",
									 -- x"8F8E9092", x"94939395", x"989A9B9B", x"9B9DA0A2", x"A2A5A8A8", x"A6A6A9AC", x"ACADAFB0", x"B2B1B0AF",
									 -- x"B0B1B1B0", x"B0B1B3B5", x"B3B7BABA", x"BCC0C3C3", x"C1C2C3C3", x"C5C7C8C7", x"C5C6C6C7", x"C7C7C6C6",
									 -- x"C3C4C4C5", x"C5C5C6C7", x"C8C7C4C1", x"C2C4C4C2", x"C3C1C0BF", x"C0BFBEBC", x"BDBDBCBD", x"BDBDBCBC",
									 -- x"BBB9B7B5", x"B4B3B2B2", x"B5B5B5B6", x"B8B8B7B5", x"BCB8B7BB", x"BDBDBEC1", x"BDBDBEBF", x"BFBFC0C0",
									 -- x"C2C3C3C1", x"C1C3C3C2", x"C3C2C1C1", x"C2C2C2C2", x"C0C1C2C2", x"C1C1C1C1", x"BEBEBEBC", x"BCBDBDBB",
									 -- x"BBBAB8B8", x"B9B9B9B9", x"B7B7B4B2", x"B5B5B5B8", x"B7B8B9BA", x"BABAB9B8", x"BCBAB7B5", x"B4B5B5B6",
									 -- x"B6B5B5B4", x"B4B3B3B3", x"B4B5B5B4", x"B3B3B3B3", x"B0AFAFB0", x"B1B1B0AF", x"B3B3B3B4", x"B4B4B4B4",
									 -- x"B8BBBAB5", x"B6BBB9B3", x"B6B4B2B1", x"B1B1B1B1", x"B1B3B5B6", x"B7B8B7B7", x"B5B7B2AE", x"AFAEABAB",
									 -- x"ACABAAAA", x"A9A8A7A6", x"A7A6A5A3", x"A1A0A0A1", x"9E9C9C9D", x"9D9C9C9C", x"969B9A94", x"93969692",
									 -- x"94979A9A", x"98969798", x"989A9997", x"999C9B97", x"95969898", x"97969595", x"94989C9A", x"98999DA0",
									 -- x"A2A7ABAC", x"AEB1B0AC", x"ACA9A6A5", x"A6A6A5A5", x"A5A4A4A5", x"A3A1A1A3", x"A2A6A7A2", x"A1A4A4A0",
									 -- x"A7AAAAA8", x"A7A9A9A8", x"A0A2A09C", x"9C9E9B96", x"91929496", x"94908E8F", x"948F8E87", x"888E8B8C",
									 -- x"87878686", x"85858586", x"85878682", x"81828281", x"7F808182", x"82817F7D", x"7C7C7C7B", x"7A7A7B7D",
									 -- x"76747577", x"777A7A74", x"7A7B7C7D", x"7D7D7C7B", x"7C7F7F7E", x"7F83837F", x"84808180", x"7A787979",
									 -- x"7D7A7C77", x"7374747C", x"79777473", x"74737270", x"6B6F7475", x"73717071", x"6D6D6E6F", x"6D6C6F74",
									 -- x"6E727779", x"79787879", x"7A7B7C7E", x"7D7B7D80", x"80818080", x"83888A8C", x"91919897", x"96979396",
									 -- x"999A9896", x"999E9F9C", x"9C9B9B9D", x"9E9D9B9B", x"969A9E9E", x"9C9A9C9E", x"9A969599", x"99949396",
									 -- x"9794908F", x"91949594", x"9692979E", x"9D9A9896", x"99989797", x"96969695", x"9D9D9D9E", x"9F9F9FA0",
									 -- x"9F9C9B9C", x"9E9EA0A2", x"A3A19FA0", x"A2A3A3A2", x"A5A5A6A7", x"A6A6A8AA", x"ACACACAD", x"AFB0B0AF",
									 -- x"B2B2AEB3", x"B5B2B4B2", x"B4B2B0B0", x"B0B0AEAD", x"AFAFB0B2", x"B2B3B3B3", x"B8B4B0B0", x"B3B6B4B1",
									 -- x"8D8D8F92", x"93949699", x"9B9C9C9C", x"9C9D9FA1", x"A2A5A7A7", x"A7A7A9AC", x"ACADAEAF", x"B0B1B1B0",
									 -- x"AEAFB0B1", x"B1B2B5B8", x"B4B7B9BA", x"BBBEC1C1", x"C1C3C4C3", x"C3C5C7C8", x"C5C6C6C6", x"C6C5C5C4",
									 -- x"C4C4C4C4", x"C4C5C5C6", x"C6C6C4C2", x"C2C4C4C2", x"C3C2C1C1", x"C1C0BFBE", x"BEBEBEBF", x"BFBEBDBC",
									 -- x"B9B7B5B3", x"B2B1B0B0", x"B2B3B4B5", x"B7B8B8B7", x"BCBAB9BB", x"BCBDBEBF", x"BEBFBFC0", x"C0C1C1C2",
									 -- x"C2C4C3C1", x"C1C3C3C1", x"C1C0BFBF", x"C0C0C0C0", x"BEBFC0C0", x"C0BFC0C0", x"C0C0BFBC", x"BCBDBCBB",
									 -- x"B9B8B7B6", x"B7B8B7B7", x"B5B6B4B4", x"B6B6B5B7", x"B6B6B7B8", x"B9B8B8B8", x"B9B7B5B4", x"B4B5B5B5",
									 -- x"B5B4B3B2", x"B2B2B3B3", x"B3B3B3B2", x"B1B1B1B1", x"B1B1B0B1", x"B1B1B0AF", x"AFB0B1B1", x"B2B3B3B3",
									 -- x"B7B8B8B7", x"B6B6B5B4", x"B4B3B1B0", x"AFB0AFAF", x"B1B2B4B5", x"B6B6B6B6", x"B4B6B2AE", x"AFAEABAA",
									 -- x"ABAAAAA9", x"A9A8A7A6", x"A7A6A5A3", x"A2A1A1A1", x"A19E9C9D", x"9C9B9A9B", x"979A9996", x"94969694",
									 -- x"96999C9D", x"9B999A9A", x"98989898", x"9A9C9B99", x"989A9B9B", x"9A999898", x"9A9A9A9B", x"9FA2A3A1",
									 -- x"A3A8ABAC", x"AFB2B3B0", x"AFAEACAB", x"ABABABAB", x"ABAAAAAB", x"AAA6A4A4", x"A6A8A7A3", x"A2A5A6A4",
									 -- x"A5A8A9A9", x"A9ABABA9", x"A5A4A3A2", x"A19E9C9A", x"97969696", x"94919192", x"908D8E89", x"898E8A8B",
									 -- x"88888787", x"86868788", x"88888784", x"83838280", x"7E7E7F7F", x"7F808182", x"7B7B7B79", x"7878797B",
									 -- x"7A777878", x"787C7E7A", x"7778797B", x"7C7C7C7C", x"7A7D7E7E", x"8083817C", x"817E7F7F", x"7B797A79",
									 -- x"78767A78", x"76757276", x"79787674", x"73737476", x"74727070", x"7272716F", x"6D6D6D6C", x"6A696D71",
									 -- x"6F727576", x"76767676", x"77787A7D", x"7D7B7979", x"7F818081", x"8687878A", x"8C8C9393", x"93959397",
									 -- x"92959695", x"979B9A96", x"9997989C", x"9F9F9E9D", x"9B9C9D9C", x"9A979696", x"96939395", x"95939396",
									 -- x"9493918F", x"8E8E9092", x"94939799", x"98999995", x"97959394", x"95969493", x"9B9B9B9B", x"9C9C9D9E",
									 -- x"9A999999", x"9A9C9E9F", x"A4A3A2A2", x"A2A19F9F", x"A3A4A5A6", x"A7A6A6A7", x"ACADADAC", x"ABAAA9A9",
									 -- x"AEAFADB3", x"B5B2B4B2", x"AFAFAFAF", x"AFAFAFB0", x"AFAFAFAF", x"B1B1B2B2", x"B6B4B2B1", x"B3B4B4B4",
									 -- x"8F8F9192", x"9293969B", x"9E9D9D9D", x"9E9F9F9F", x"A2A3A5A6", x"A6A8A9AA", x"ACACADAE", x"AFB0B2B2",
									 -- x"B2B2B3B2", x"B1B2B4B5", x"B5B7B9B9", x"BABDBFC0", x"C1C4C5C3", x"C1C3C6C8", x"C6C6C5C5", x"C4C4C3C2",
									 -- x"C5C3C2C2", x"C3C4C4C4", x"C5C5C4C3", x"C3C4C4C3", x"C1C2C2C1", x"C0BFBEBE", x"BDBEBFBF", x"BEBDBCBC",
									 -- x"B8B7B4B2", x"B1B1B1B0", x"AFB0B3B5", x"B6B7B8B9", x"BABBBABA", x"BBBDBDBB", x"BFBFC0C0", x"C1C1C2C2",
									 -- x"C2C3C3C1", x"C1C2C1C0", x"BFBFBEBF", x"BFBFBFBE", x"BEBFC0C0", x"C0C0C1C1", x"C1C1BFBC", x"BCBDBCBA",
									 -- x"B8B7B6B6", x"B6B6B6B5", x"B3B6B5B5", x"B7B6B3B5", x"B3B3B4B5", x"B5B6B6B7", x"B6B5B4B3", x"B4B4B4B4",
									 -- x"B4B3B1B0", x"B0B1B2B2", x"B0B1B1B0", x"AFAEAEAE", x"B1B1B0B0", x"B0AFAEAD", x"AEAEAFB0", x"B1B1B2B2",
									 -- x"B2B1B3B5", x"B3AEAEB2", x"B1B0AFAE", x"AEAEAEAE", x"B0B1B2B4", x"B5B5B5B5", x"B3B5B1AE", x"AEADAAA9",
									 -- x"AAA9A9A9", x"A9A8A6A5", x"A6A6A5A4", x"A3A2A1A1", x"A3A09D9D", x"9C9B9B9C", x"99999897", x"96959596",
									 -- x"989B9E9F", x"9E9C9C9C", x"9C9A9A9B", x"9B999898", x"9B9B9C9C", x"9B9A9A9A", x"9C9B9B9E", x"A3A7A6A3",
									 -- x"A5A9ACAD", x"B0B5B6B4", x"B1B1B0AF", x"AEAEAFB0", x"AFADADAE", x"AEAAA7A5", x"A9A8A5A4", x"A4A5A7A8",
									 -- x"A5A8AAAA", x"ABACABA9", x"A5A2A1A4", x"A39D9B9D", x"9A979595", x"94929191", x"8D8D908C", x"8B8D898A",
									 -- x"8B8A8A89", x"88888889", x"8A8A8885", x"8584827F", x"7D7D7E7E", x"7E7F8081", x"7B7A7978", x"77777879",
									 -- x"75757878", x"77787975", x"7A7A7979", x"78777676", x"78797A7A", x"7D81807C", x"807D7D7E", x"78757574",
									 -- x"74717675", x"75746E70", x"72757878", x"76737170", x"74747370", x"6C6C6E71", x"70706F6E", x"6C6B6E72",
									 -- x"71717171", x"72727272", x"7575787D", x"7E7C7876", x"7B7E7C7F", x"87848186", x"8989908F", x"90949296",
									 -- x"90939594", x"94979795", x"9896979C", x"A0A1A09F", x"A09E9D9B", x"99969492", x"96959492", x"91909091",
									 -- x"9091918F", x"8B8B8F92", x"92959897", x"95999B96", x"94918F90", x"94959391", x"99999999", x"9A9A9B9B",
									 -- x"989A9A97", x"989C9D9C", x"A0A2A3A2", x"A2A1A1A0", x"A1A2A4A6", x"A7A7A5A3", x"A8AAACAC", x"ABABACAE",
									 -- x"ABAEADB2", x"B3AFB2B0", x"ADAEAFAE", x"ADADAEB0", x"AFADADAD", x"AFB0B0AF", x"B1B1B2B2", x"B1B2B3B5",
									 -- x"94949494", x"91919499", x"9E9D9C9D", x"9FA0A09F", x"A1A1A2A4", x"A6A7A8A8", x"ABACADAE", x"AFB0B1B2",
									 -- x"B3B4B4B4", x"B2B2B3B4", x"B5B6B7B8", x"BABDBFC0", x"C2C4C4C2", x"C1C3C4C5", x"C5C5C4C4", x"C3C3C2C2",
									 -- x"C5C2C0C0", x"C2C4C4C3", x"C4C4C4C4", x"C4C4C3C2", x"BFC0C1C0", x"BEBDBDBD", x"BBBDBFBF", x"BDBBBABA",
									 -- x"B8B6B3B2", x"B1B1B1B1", x"ADAFB2B4", x"B5B6B9BA", x"B8BBBBB9", x"BABDBCB9", x"BEBEBEBF", x"C0C1C1C1",
									 -- x"C1C2C1C1", x"C0C0C0BF", x"C0C0BFBF", x"C0C0BFBE", x"BEBFC0C0", x"C0C0C1C1", x"BFBFBEBC", x"BBBCBBB9",
									 -- x"B8B7B7B7", x"B7B6B5B5", x"B3B6B5B5", x"B6B4B1B3", x"B1B1B1B2", x"B3B4B5B6", x"B6B5B4B4", x"B4B3B2B2",
									 -- x"B2B2B1B0", x"B0AFAFB0", x"ADAEAEAE", x"ADADADAD", x"AFAFAEAE", x"AEAEADAC", x"AFB0B0B0", x"B1B1B0B0",
									 -- x"AEAEAFB1", x"B0ADADAF", x"B0AFAEAD", x"AEAEAEAE", x"B0B1B2B3", x"B4B4B4B4", x"B1B4B1AD", x"AEADA9A8",
									 -- x"A9A9A8A9", x"A9A8A6A5", x"A5A5A4A4", x"A4A4A3A3", x"A4A19E9D", x"9D9C9D9F", x"99979798", x"97949497",
									 -- x"999C9FA0", x"9E9C9B9B", x"9D9B9A9C", x"9C99989A", x"9D9E9E9E", x"9E9D9D9D", x"9B9FA1A2", x"A4A7A9A9",
									 -- x"A8ACAFB0", x"B3B6B7B5", x"B3B4B3B2", x"B0B0B1B3", x"B1AEADAF", x"B0AEABA9", x"AEAAA7A8", x"A8A7A9AC",
									 -- x"AAAAABAC", x"ACABA9A7", x"A3A0A0A2", x"A09D9C9F", x"99979697", x"97949190", x"8F8F938F", x"8C8D898B",
									 -- x"8E8D8B8A", x"8A898988", x"8B898684", x"8484817E", x"7D7D7D7F", x"807F7D7B", x"7B7A7977", x"77777778",
									 -- x"78797B7B", x"77797B78", x"7C7B7977", x"76747373", x"77767574", x"787E8180", x"807C7C7C", x"78757573",
									 -- x"736F7270", x"70706C6F", x"70737678", x"76726F6D", x"6F717270", x"6B696B6D", x"7171716F", x"6E6E7072",
									 -- x"71706E6D", x"6E6F7070", x"7373777A", x"7B797777", x"797B787C", x"84827E85", x"88878C8C", x"8D908F92",
									 -- x"9092928F", x"8E919496", x"9997979B", x"9F9F9D9B", x"9E9D9B99", x"97949392", x"95969591", x"8F8F8F8D",
									 -- x"8B8D8E8D", x"8B8B8F93", x"90929595", x"94979A97", x"928F8E8E", x"90939393", x"96979899", x"9A9B9B9A",
									 -- x"979B9B97", x"979C9D9A", x"9DA0A1A1", x"A0A1A2A2", x"A0A1A3A4", x"A6A7A5A2", x"A4A5A8AA", x"ADAFB1B2",
									 -- x"ABAFAEB2", x"B0ABAEAE", x"AEAFAFAE", x"ACABABAC", x"ADACABAD", x"AFB0AEAD", x"ADAEAFAF", x"AFB0B1B3",
									 -- x"95959595", x"92919599", x"9D9C9C9D", x"9FA1A1A1", x"A2A2A2A4", x"A6A8A8A8", x"AAACADAF", x"AFAFB0B1",
									 -- x"B0B2B3B4", x"B3B3B5B6", x"B4B4B6B8", x"BBBEC0C2", x"C2C2C2C2", x"C3C4C3C0", x"C3C3C3C3", x"C3C3C3C3",
									 -- x"C3C0BEBF", x"C1C3C4C3", x"C4C4C4C4", x"C3C2C1C1", x"BEC0C1C0", x"BEBCBCBD", x"BCBDBEBE", x"BDBBB9B8",
									 -- x"B5B3B0AF", x"AFAFB0B0", x"AEB0B2B4", x"B4B5B7B9", x"B8BCBDBB", x"BBBDBDBA", x"BFBEBEBF", x"C0C1C0C0",
									 -- x"C1C1C1C1", x"C1C0C0BF", x"C1C0BFBF", x"BFBEBEBD", x"BCBDBEBE", x"BDBDBDBE", x"BCBDBCBA", x"BABAB8B5",
									 -- x"B7B7B7B7", x"B6B5B4B4", x"B3B6B5B3", x"B3B1AEB1", x"B0B0B0B1", x"B2B3B5B6", x"B5B5B4B4", x"B3B3B2B1",
									 -- x"B1B1B2B1", x"B0AEADAC", x"ABACACAC", x"ABACADAE", x"ADADADAD", x"AEAEADAC", x"AFAFAFB0", x"B0B0AFAF",
									 -- x"ADAEAFAE", x"B0B1B0AE", x"AFAEADAD", x"AEAEAFAF", x"B0B0B1B2", x"B3B3B3B3", x"B0B3B0AC", x"ADACA8A8",
									 -- x"A9A9A9A9", x"A9A8A7A5", x"A4A4A3A4", x"A5A5A4A4", x"A4A19E9E", x"9D9C9D9E", x"9A979799", x"98949598",
									 -- x"9B9D9FA0", x"9F9D9C9B", x"9C9A9A9D", x"9E9B9B9E", x"A1A1A2A2", x"A3A3A2A1", x"A0A3A6A6", x"A7AAACAD",
									 -- x"ABAEB1B3", x"B5B7B7B6", x"B7B7B7B6", x"B4B3B4B5", x"B6B2B0B1", x"B2B2B0B0", x"B2ADABAD", x"AEACACAF",
									 -- x"AEADADAD", x"ADABA9A8", x"A4A3A2A0", x"A0A0A1A1", x"9B99989A", x"9A989595", x"92919592", x"8F8F8C90",
									 -- x"8F8D8C8B", x"8B8B8A89", x"8C898584", x"84838280", x"807D7C7D", x"80807B76", x"7A797876", x"76757575",
									 -- x"7A797876", x"72767D7D", x"78777676", x"75767676", x"75757373", x"767B7F80", x"7D797A7B", x"79787978",
									 -- x"716E716F", x"6D6F6D73", x"76737170", x"70727373", x"726D6A6B", x"6E6F6B67", x"6C6D6E6E", x"6D6E6E6F",
									 -- x"716F6E6D", x"6E707171", x"71727475", x"74727377", x"7C7D7A7B", x"807F7F86", x"85848989", x"8A8D8B8E",
									 -- x"8E8F8E8B", x"8A8C9093", x"98969699", x"9C9A9796", x"98989795", x"92909091", x"8F909190", x"90908F8D",
									 -- x"8889898A", x"8A8C8E90", x"8E8C9094", x"92919292", x"90908E8D", x"8D909396", x"92959898", x"9A9B9B98",
									 -- x"94989996", x"969A9B98", x"9EA0A19E", x"9D9EA0A0", x"A0A1A2A2", x"A4A7A5A2", x"A5A4A4A6", x"AAACABAA",
									 -- x"ACAFADB0", x"ADA8ACAD", x"B0AFAEAD", x"ACABA9A8", x"AAAAABAD", x"AFAFAEAC", x"AEADADAE", x"AFB1B1B1",
									 -- x"92929495", x"9595999D", x"9C9C9D9E", x"A0A1A2A2", x"A4A4A4A5", x"A7A9A9A9", x"A8AAADAE", x"AEAEAFB0",
									 -- x"B0B2B3B4", x"B3B3B3B4", x"B5B4B5B8", x"BBBDC0C2", x"C2C2C1C1", x"C4C5C2BE", x"C1C1C1C1", x"C1C2C2C3",
									 -- x"C0BFBEBF", x"C0C2C3C2", x"C3C3C3C3", x"C2C0C0C1", x"C0C0C0BF", x"BEBEBEBE", x"BEBDBDBD", x"BDBBB9B7",
									 -- x"B3B1AFAD", x"AEAEAFB0", x"AFB0B1B2", x"B3B4B5B6", x"B9BBBCBC", x"BCBDBEBD", x"C0BFBEBF", x"C0C0C0BF",
									 -- x"C1C0C0C2", x"C2C0BFC0", x"C0BEBCBB", x"BABABAB9", x"BBBCBCBC", x"BCBBBBBC", x"BABBBAB8", x"B7B7B5B2",
									 -- x"B5B5B5B4", x"B3B2B2B2", x"B2B5B3B1", x"B0ADABAE", x"AFAFAFB0", x"B1B2B4B5", x"B2B1B1B1", x"B2B2B2B1",
									 -- x"B0B1B1B1", x"B0ADAAA9", x"AAAAAAAA", x"AAABAEAF", x"ADADADAE", x"AFAFAFAE", x"ACACADAD", x"AEAEAEAE",
									 -- x"ABADACAB", x"ADB0AFAB", x"AFADACAC", x"ACAEAFAF", x"B0B0B1B1", x"B2B2B2B2", x"B0B2AEAB", x"ACABA7A7",
									 -- x"A9A9A9AA", x"AAA9A8A6", x"A5A4A4A4", x"A6A6A5A3", x"A3A19E9E", x"9D9B9A9B", x"9A98989A", x"99969799",
									 -- x"9D9FA0A1", x"A09E9D9D", x"9E9E9E9F", x"9E9C9B9D", x"A1A1A2A4", x"A5A5A4A3", x"A4A3A3A4", x"A9ADADAA",
									 -- x"ADB0B3B6", x"B8B9B9B8", x"BABAB9B8", x"B7B6B6B7", x"BBB8B4B4", x"B4B3B3B4", x"B2AEADAE", x"AFADACAD",
									 -- x"B0AEADAE", x"AFADABAA", x"A7A6A3A0", x"A0A2A1A0", x"9E9B9998", x"9898999A", x"96949794", x"92929095",
									 -- x"8F8D8B8B", x"8C8D8C8B", x"8C898686", x"85848382", x"827E7A7B", x"7E7F7C78", x"78777575", x"74737271",
									 -- x"70717575", x"73767977", x"76757574", x"74757576", x"72747575", x"76777879", x"7A767779", x"77767775",
									 -- x"6E6C706F", x"6E6F6E73", x"706E6C6C", x"6F717272", x"716E6A69", x"6B6C6C6A", x"686A6C6C", x"6C6D6D6D",
									 -- x"6F6F6E6E", x"6F707172", x"72737573", x"706E7176", x"7C7B7C7B", x"7A7C8082", x"83828889", x"8B8E8B8D",
									 -- x"8A8C8D8D", x"8C8D8F91", x"9896979A", x"9B999695", x"95959593", x"908E8F90", x"8E8C8C8D", x"8E8D8A87",
									 -- x"8A8A8A8A", x"8C8E8E8F", x"908B8E93", x"928E8E8D", x"908F8E8C", x"8B8D9296", x"8F939696", x"979A9996",
									 -- x"91969897", x"979A9B9A", x"9A9D9D9B", x"9B9EA09F", x"9FA1A2A1", x"A2A5A5A3", x"A6A4A2A4", x"A7A9A7A4",
									 -- x"AAADABAE", x"ACA8ACAC", x"AEADACAC", x"ADACA9A7", x"A8A9ABAD", x"AEAEADAD", x"B1AEADAE", x"B0B2B1B0",
									 -- x"90909296", x"98999B9E", x"9D9E9FA0", x"A0A0A1A2", x"A4A4A5A6", x"A6A7A8A9", x"A6A8AAAB", x"ABACAEB0",
									 -- x"B0B2B4B4", x"B2B1B1B1", x"B7B5B4B7", x"BABBBDBF", x"C1C1C1C1", x"C2C3C2BF", x"BFBFBFBF", x"BFC0C1C2",
									 -- x"BFBFBFBF", x"C0C0C1C1", x"C2C1C2C2", x"C1BFBFC2", x"C1C0BFBE", x"BEBEBEBE", x"BFBDBBBB", x"BCBBB8B6",
									 -- x"B2B0AEAC", x"ADAEAFB0", x"B0AFAFB0", x"B1B2B3B3", x"B7B7B9BB", x"BBBBBCBE", x"C0BFBDBE", x"BFBFBEBC",
									 -- x"BEBDBDC0", x"C0BEBDBE", x"BEBCB9B7", x"B6B6B5B5", x"B8B9BABA", x"BABABABA", x"B8B8B7B5", x"B5B6B5B3",
									 -- x"B4B4B4B2", x"B0AFB0B1", x"B0B3B2AF", x"AEABA9AC", x"ABABACAD", x"AEAFB0B0", x"AFAFAEAE", x"AFB0B0AF",
									 -- x"AFAFB0AF", x"AEACA9A8", x"AAAAA9A8", x"A8AAADAF", x"ADADADAE", x"AFAFAFAF", x"AAABABAC", x"ADADADAD",
									 -- x"AAA8A8A8", x"A9A9A9AA", x"ADABAAA9", x"AAACAEAF", x"AFAFB0B0", x"B0B1B1B1", x"AFB1ADAA", x"ABAAA7A7",
									 -- x"A9AAAAAB", x"ACABA9A7", x"A7A6A5A5", x"A6A6A4A2", x"A2A09FA0", x"9F9D9B9B", x"9B9B9B9B", x"9A999A9B",
									 -- x"9E9E9FA0", x"A09F9F9F", x"A0A2A29F", x"9D9D9C9C", x"9FA0A2A5", x"A6A7A5A3", x"A3A2A2A2", x"A6ABACAB",
									 -- x"AFB0B3B7", x"BABCBDBD", x"BDBCBCBB", x"BCBBBBBA", x"BEBBB8B6", x"B5B4B5B7", x"B3B0AEAD", x"AEAEADAC",
									 -- x"B1AFAFB1", x"B1AFABAA", x"A9A4A1A2", x"A4A29F9F", x"9F9C9A9A", x"99989A9D", x"9B979997", x"94949196",
									 -- x"918F8D8C", x"8D8E8D8B", x"8A888888", x"86838182", x"817F7C7C", x"7C7C7B79", x"76757575", x"7473706E",
									 -- x"6E70777A", x"797A7975", x"76767573", x"72717170", x"70737576", x"74727476", x"78747678", x"7573726E",
									 -- x"6F6B6D6C", x"6B6D6A6E", x"67696B6D", x"6E6E6C6B", x"6D6F6F6B", x"6665696E", x"67696B6A", x"6B6D6D6C",
									 -- x"6A6C6E6E", x"6E6E6F70", x"72737473", x"716F7175", x"77767D7C", x"747A817D", x"80808788", x"8B8E898B",
									 -- x"87898C8F", x"8F8F8F90", x"9696989A", x"99969494", x"93939291", x"908F8F8E", x"918B888B", x"8C898482",
									 -- x"89898A8A", x"8B8C8D8D", x"918D8E91", x"90908F8B", x"8F8E8C8B", x"8B8C8F92", x"90939594", x"95989794",
									 -- x"92949798", x"9797999A", x"97999A99", x"9B9FA09D", x"9CA0A2A0", x"A0A4A4A2", x"A4A3A2A4", x"A6A7A6A4",
									 -- x"A7AAA8AC", x"ABA7ABAA", x"A9AAABAC", x"ACABA9A7", x"A8AAABAC", x"ABABACAE", x"B3B0AEAE", x"B0B1B1B0",
									 -- x"91919397", x"999A9B9D", x"9FA0A2A1", x"A0A0A1A2", x"A2A3A4A5", x"A5A5A6A7", x"A5A6A8A8", x"A9AAAEB1",
									 -- x"ACAFB1B3", x"B3B2B3B3", x"B9B6B4B7", x"B9B9BABC", x"C0C2C2C0", x"C0C2C2C1", x"BEBEBDBD", x"BEBFC0C0",
									 -- x"BEBFC0BF", x"BFBFBFC0", x"C1C0C0C2", x"C1BFC0C3", x"C1BFBDBC", x"BDBDBDBD", x"BEBBB9B9", x"BABAB7B4",
									 -- x"AFADABA9", x"AAABADAD", x"B0AFAEAE", x"B0B1B1B0", x"B5B4B5B9", x"BAB8BABE", x"BFBDBCBC", x"BDBDBCBA",
									 -- x"BAB9BABD", x"BDBBBABC", x"BEBBB8B5", x"B4B3B3B3", x"B4B5B6B7", x"B7B7B7B8", x"B6B6B4B3", x"B4B6B8B7",
									 -- x"B4B4B3B1", x"AFAFB0B1", x"ADB1B1AF", x"AEAAA8AA", x"A7A8A8A9", x"AAABACAC", x"AEADACAC", x"ACACACAC",
									 -- x"AEAEAEAD", x"ACAAA9A8", x"ABAAA8A7", x"A7A9ACAF", x"ACACACAD", x"AEAEAEAD", x"ACACACAC", x"ACACACAB",
									 -- x"ABA7A6AA", x"A8A3A5AB", x"ACAAA8A7", x"A8AAADAE", x"AEAEAFAF", x"AFAFB0B0", x"AFB1ADA9", x"AAA9A7A7",
									 -- x"AAAAABAC", x"ACACAAA8", x"A8A7A5A5", x"A6A5A3A0", x"A2A0A1A2", x"A2A09E9E", x"9C9D9D9B", x"9B9B9C9C",
									 -- x"9D9D9E9F", x"9FA0A0A0", x"9B9FA19F", x"9EA1A2A0", x"A0A1A3A7", x"A9A9A7A5", x"A0A4A7A5", x"A4A7ACB0",
									 -- x"AFB0B3B7", x"BBBEC0C2", x"C2C1C0C0", x"C1C2C1BF", x"BFBDBBB9", x"B8B6B8BB", x"B7B5B2AF", x"B0B1B0AE",
									 -- x"B2B0B0B3", x"B3AFABA9", x"ABA29FA6", x"A9A39FA1", x"9F9F9F9F", x"9D9B9C9E", x"9F9A9C98", x"96949094",
									 -- x"94928F8E", x"8E8D8B8A", x"87878889", x"86817F7F", x"7F7F807F", x"7D7B7877", x"76767576", x"7573706E",
									 -- x"73717171", x"6F737775", x"74747372", x"716F6F6E", x"6F727473", x"706F7377", x"7673767B", x"79767470",
									 -- x"736B6A66", x"66686568", x"6A6B6C6C", x"6A6A6B6D", x"6D6D6C6A", x"67666667", x"66696968", x"696B6C6B",
									 -- x"65686C6C", x"6B6B6B6C", x"6E6E7072", x"71707173", x"72737F7F", x"747C867D", x"7C7C8385", x"87898484",
									 -- x"8485888B", x"8D8E8F90", x"93949697", x"95919090", x"908F8D8E", x"8F8F8E8C", x"91888489", x"8C898584",
									 -- x"84858687", x"8788898A", x"8D8C8C8C", x"8D929189", x"8E8C8A8A", x"8B8C8D8D", x"92959593", x"93979794",
									 -- x"91929496", x"95929395", x"989A9A98", x"9A9D9C97", x"9A9FA2A0", x"A0A2A3A1", x"A3A3A3A3", x"A4A4A3A3",
									 -- x"A6A8A7AC", x"ABA7A9A7", x"A6A8ABAC", x"ABA9A8A7", x"A8AAABAA", x"A8A8ABAE", x"B2B0AEAD", x"AEAFAFAF",
									 -- x"9094999A", x"99999B9E", x"9E9E9F9F", x"9FA1A2A3", x"A3A1A3A6", x"A9A8A8A8", x"A8A7A6A7", x"ABAFAEAC",
									 -- x"B0AEAEB0", x"B2B1B2B4", x"B5B5B6B8", x"BABCBDBD", x"BEC0C2C3", x"C3C1C0BF", x"BDBDBDBE", x"BFBFC0C1",
									 -- x"C2BFBDBC", x"BDBEBFC0", x"C0BFC0C2", x"C2BFBDBD", x"C0BEBCBC", x"BDBEBEBE", x"BCBCBAB9", x"B8B7B5B4",
									 -- x"ADACAAAB", x"ACADACAB", x"ABADAFAF", x"AEAEB1B3", x"B2B1B3B7", x"B9B8B7B9", x"BFBEBAB7", x"B7B9B8B5",
									 -- x"B8B7B7B8", x"B9B9B8B7", x"B7B7B7B5", x"B3B1AFAF", x"ACAEB0B2", x"B3B3B3B3", x"B0B0B0B1", x"B2B2B2B1",
									 -- x"B4B2B0AF", x"AFAFAFAF", x"B1AFACAB", x"ABABA9A7", x"A6A7A8A8", x"A8A8A8A9", x"ABADADAA", x"A9ABADAD",
									 -- x"ABACADAD", x"ACABABAB", x"A6A8A8A6", x"A7AAACAC", x"ABA9AAAE", x"B0AEADAF", x"ADAFADAA", x"ABAEACA8",
									 -- x"A9A8A7A5", x"A5A5A6A7", x"A7A6A5A5", x"A6A8AAAC", x"AEAFB0AE", x"ADAEAFAE", x"AEB0B0AD", x"AAAAAAAA",
									 -- x"AAA9A9AB", x"ACAAA8A7", x"A5A5A5A5", x"A6A6A4A3", x"A4A2A1A0", x"A0A09F9F", x"9B9B9C9D", x"9D9D9C9B",
									 -- x"9F9E9E9F", x"9E9EA0A3", x"9E9FA09F", x"9D9EA2A5", x"A3A1A5A9", x"A6A6A9AA", x"A9A8A7A6", x"A6A9ACAF",
									 -- x"B0B4B7B7", x"B9BCC1C3", x"C2C0BFC0", x"C3C5C4C3", x"C3C0BDBC", x"BDBDBCBA", x"B6B6B5B2", x"AFAFB2B5",
									 -- x"B3B3B1AF", x"AFB1AFAB", x"AAA8A8A8", x"A7A3A2A3", x"A4A2A0A0", x"A1A2A1A0", x"9D9C9C9C", x"9B9A9694",
									 -- x"95939394", x"918C8B8E", x"8D8B8986", x"85848382", x"7C7D7D7C", x"7E7F7C77", x"76757472", x"70706F6D",
									 -- x"73727171", x"72727271", x"71716D6A", x"6B6F6E6A", x"6C6E7071", x"6F6E7175", x"6F757A78", x"74706E6C",
									 -- x"6D696668", x"6A696767", x"6B696C6E", x"6B6C6E6C", x"6F6C6A6B", x"69656568", x"696A6D6C", x"67686A68",
									 -- x"67706D68", x"6D6B676C", x"6B68676B", x"6F706F6F", x"7274777A", x"7B7C7F83", x"7F808589", x"87828288",
									 -- x"8C88878B", x"8B898D94", x"8F919190", x"8F8F8E8C", x"8C90928E", x"8988898A", x"898A8883", x"82858889",
									 -- x"86878786", x"85848586", x"878A8B8A", x"8B8F8E8B", x"8A88878C", x"93918D8F", x"8D909292", x"94959592",
									 -- x"9091908E", x"8F929392", x"95979A9A", x"9998999B", x"9F9F9E9E", x"9FA0A2A3", x"A0A1A2A3", x"A4A5A5A5",
									 -- x"A4A5A6A7", x"A9ABA8A4", x"A2A6AAA9", x"A6A4A6A9", x"ACA9ABAA", x"A6ABB1AE", x"ADADAEB1", x"B2B1AEAA",
									 -- x"93959798", x"999A9C9E", x"9FA0A0A1", x"A1A2A4A5", x"A3A2A3A6", x"A8A7A7A7", x"A9A8A7A7", x"A9ACADAE",
									 -- x"AEAFB1B3", x"B2B1B2B4", x"B5B5B5B7", x"B9BCBDBD", x"BEC0C1C2", x"C2C0BFBE", x"BDBDBEBE", x"BEBEBEBE",
									 -- x"BEBCBAB9", x"BABCBDBD", x"BFBFC0C2", x"C2BFBEBE", x"BEBDBCBD", x"BEBEBEBD", x"BCBBB9B8", x"B6B4B2B1",
									 -- x"ACABAAAA", x"AAABABAB", x"A7A8AAAC", x"AEAFAFAF", x"B4B3B4B5", x"B5B4B6B9", x"BABAB8B6", x"B5B8B8B7",
									 -- x"B6B6B5B6", x"B7B7B6B6", x"B5B5B5B4", x"B2B0AEAD", x"A8A8A9AC", x"AFB1B1B0", x"AEAEAFAF", x"B0B0B0AF",
									 -- x"B1B0AFAF", x"AFAFAFAF", x"ADABAAA9", x"AAAAA8A6", x"A4A3A4A6", x"A8AAAAA9", x"A7AAADAC", x"ABACABA9",
									 -- x"A9A9AAAA", x"AAA9A9A9", x"A7A9A9A8", x"A8ABADAC", x"ABAAABAE", x"AFAEAEAE", x"ACADACA9", x"AAADABA7",
									 -- x"A8A7A6A5", x"A5A6A6A7", x"A9A9A8A7", x"A7A8AAAB", x"A9ABADAD", x"ADAEAFAE", x"ADAEADAA", x"A8A9A8A7",
									 -- x"A9AAABAB", x"AAA8A7A7", x"A7A7A6A6", x"A6A6A6A5", x"A6A4A2A0", x"9F9E9D9C", x"9C9D9F9F", x"9E9E9E9F",
									 -- x"A09F9FA0", x"9F9EA0A2", x"A1A19F9E", x"9D9FA0A2", x"A4A2A5A8", x"A6A6A8A8", x"A7A8A8A9", x"A9ABACAE",
									 -- x"B3B5B8B9", x"BCC1C4C5", x"C5C4C3C3", x"C2C2C1C1", x"C4C1BEBE", x"C0C0BDBA", x"BAB9B7B5", x"B2B2B3B4",
									 -- x"B4B5B3B2", x"B2B2AFAB", x"ACAAA9A9", x"A8A6A6A8", x"A4A4A4A4", x"A3A2A3A3", x"A5A3A09E", x"9D9B9997",
									 -- x"96969797", x"95918F90", x"8C8A8887", x"86858383", x"83807E7F", x"7D797676", x"7373716F", x"6E6D6E6E",
									 -- x"6F6F7071", x"7171706F", x"6D6E6F6E", x"6D6D6C6A", x"6C6B6C6E", x"6F6F7071", x"70737573", x"71706F6D",
									 -- x"6F6A6767", x"6767686A", x"6E6B6B6A", x"67696D6D", x"6B69696A", x"6A696A6B", x"6C6A6A68", x"65686B69",
									 -- x"6A6E6965", x"696A676A", x"6A6B6B6A", x"6C717474", x"71747779", x"7A7C7E7F", x"7C808384", x"83838483",
									 -- x"858B8D8A", x"8B919390", x"90939495", x"9595928E", x"8B8E8F8C", x"8A898988", x"87888886", x"85878887",
									 -- x"83858686", x"84848587", x"89888582", x"848A8C89", x"85888A8C", x"8C898A92", x"8C90908D", x"8A8C9195",
									 -- x"92939290", x"9091908E", x"90949798", x"98999895", x"9D9C9C9C", x"9D9E9F9F", x"A3A3A4A5", x"A5A5A5A5",
									 -- x"A3A5A6A6", x"A7A8A7A5", x"AAA6A2A1", x"A3A6A7A7", x"ACA9A8A8", x"A7A9ACAB", x"ACABACAE", x"B0B1B0AF",
									 -- x"96969697", x"999B9D9E", x"9FA0A1A1", x"A2A3A4A5", x"A5A4A5A7", x"A8A7A7A7", x"A8A9AAAA", x"A9AAABAD",
									 -- x"ACAEB1B3", x"B1AFB0B3", x"B5B4B5B6", x"B9BBBCBD", x"BEBFC0C1", x"C1BFBEBD", x"BEBEBEBD", x"BDBCBCBB",
									 -- x"BDBCBABA", x"BBBCBCBC", x"BDBCBDBF", x"BFBEBDBE", x"BBBCBDBE", x"BFBEBDBC", x"BCBBB9B7", x"B4B2AFAD",
									 -- x"AAAAA9A8", x"A8A8AAAB", x"A6A6A7AB", x"AFB1B0AD", x"B3B2B3B3", x"B3B2B5B7", x"B5B7B6B4", x"B3B4B6B7",
									 -- x"B3B3B3B4", x"B4B5B4B3", x"B1B1B2B1", x"AFACAAAA", x"A6A4A4A7", x"ABADADAB", x"ABABACAC", x"ADADADAD",
									 -- x"AFAFAEAE", x"AFAEAEAD", x"A9A8A7A8", x"A9A8A7A5", x"A6A4A3A4", x"A7A8A7A5", x"A5A8ABAB", x"ABABA9A7",
									 -- x"A8A8A8A8", x"A8A8A8A9", x"A6A7A8A7", x"A7A9ABAB", x"ABACADAD", x"AEB0AFAD", x"ABACABA9", x"AAACABA8",
									 -- x"A7A6A6A5", x"A5A5A6A7", x"A8A8A8A8", x"A8A9A9A9", x"A6AAACAC", x"ADAEADAC", x"ACACAAA8", x"A7A8A8A6",
									 -- x"A7ABADAA", x"A7A8A8A7", x"A9A8A8A6", x"A5A5A6A7", x"A6A5A2A0", x"9F9E9D9C", x"9DA0A2A1", x"9F9FA1A3",
									 -- x"A2A1A1A1", x"A09FA0A2", x"A4A29F9E", x"9FA0A1A1", x"A7A4A7AA", x"A9A9ABA9", x"A9A9AAAA", x"ABACAEB0",
									 -- x"B6B7B8BA", x"BDC2C4C3", x"C4C4C5C4", x"C3C2C2C3", x"C5C3C1C1", x"C3C2BFBB", x"BEBCBAB8", x"B7B7B6B6",
									 -- x"B4B5B5B5", x"B5B4B0AC", x"ACAAA8A8", x"A8A8A9AB", x"A5A7A8A8", x"A6A6A7A8", x"AAA8A5A3", x"A2A09E9C",
									 -- x"96989998", x"9694928F", x"8C8B8A89", x"88878584", x"857E7B7E", x"7D777578", x"6F6F6F6D", x"6C6B6C6D",
									 -- x"6D6D6E6F", x"706F6E6C", x"6D6D6E6F", x"6D6A696A", x"6A68686B", x"6F6F6D6D", x"7071716F", x"6F6F6C68",
									 -- x"67666563", x"62616265", x"69666666", x"63656968", x"69696868", x"6A6C6C6B", x"6B696867", x"666A6D69",
									 -- x"696A6969", x"6A6A6765", x"6A70726C", x"6A6F7271", x"72757777", x"797C7D7B", x"7B828480", x"81878680",
									 -- x"8484888E", x"8F8D8D8F", x"8C8D8D8E", x"90918E89", x"8E8C8885", x"86898A8A", x"87888A89", x"89898886",
									 -- x"81838686", x"84848689", x"88888886", x"888B8A86", x"84878989", x"88848790", x"8B8E908E", x"8B8B8E8F",
									 -- x"92929190", x"8F8F8D8B", x"8F939595", x"979B9A95", x"9C9C9C9C", x"9C9D9E9E", x"A2A2A2A2", x"A2A2A2A2",
									 -- x"A0A3A5A4", x"A3A4A5A5", x"A6A6A4A1", x"A0A2A6AB", x"ABA8A4A6", x"AAA9A8AB", x"ACAAA9AA", x"ADB0B1B1",
									 -- x"97979899", x"9B9C9E9F", x"9FA0A1A2", x"A2A3A4A5", x"A8A7A7A9", x"AAA8A8A9", x"A7A8AAAC", x"ACAAAAAB",
									 -- x"AEB0B1B2", x"B1B1B1B2", x"B5B5B5B6", x"B8BABBBC", x"BDBDBEBF", x"BFBFBDBC", x"BEBEBEBD", x"BCBBBABA",
									 -- x"BCBCBBBB", x"BBBCBCBC", x"BCBBBCBE", x"BEBDBCBD", x"BBBCBDBE", x"BEBDBCBB", x"BCBBB9B7", x"B4B1AEAB",
									 -- x"A8A8A8A7", x"A5A6A9AB", x"A6A6A7AA", x"AEB0AFAE", x"AEAEB0B2", x"B4B4B4B4", x"B4B4B3B2", x"B1B2B2B2",
									 -- x"B1B1B1B2", x"B2B3B2B1", x"ADADAEAD", x"AAA7A5A4", x"A4A4A5A7", x"A9AAA9A8", x"A7A8A8A9", x"AAAAACAC",
									 -- x"AEAEADAD", x"ADACAAA9", x"A8A7A7A7", x"A7A8A7A6", x"A6A5A3A4", x"A5A6A5A3", x"A6A7A7A7", x"A8A8A9A9",
									 -- x"A9A9A9A8", x"A7A7A8A9", x"A5A7A7A7", x"A7A8A9A9", x"ABAEAFAD", x"AEB0AFAC", x"ACACABAA", x"ABADACA9",
									 -- x"A7A6A5A5", x"A5A5A5A6", x"A5A5A6A7", x"A7A8A8A8", x"A8ABACAC", x"ABACABAA", x"ABAAA8A7", x"A8A9A9A7",
									 -- x"A6ABADA9", x"A7AAAAA7", x"A8A9A8A7", x"A5A4A5A6", x"A6A4A2A0", x"A0A09F9F", x"9FA0A1A1", x"A1A1A3A4",
									 -- x"A3A2A1A2", x"A2A1A1A3", x"A4A2A09F", x"A0A2A4A5", x"A8A4A6AB", x"ACADAEAC", x"AEADACAB", x"ABAEB2B5",
									 -- x"B8BABBBB", x"BDC0C1C1", x"C2C3C4C4", x"C4C4C5C5", x"C5C4C3C3", x"C3C2C0BE", x"BFBDBBBB", x"BCBCBBBA",
									 -- x"B6B6B6B6", x"B5B4B0AE", x"ACAAA9A9", x"A9A9ABAC", x"A7A9ABAB", x"ABACACAD", x"ABAAAAAA", x"AAA7A3A0",
									 -- x"999C9C98", x"9695938F", x"8E8E8D8C", x"8B898785", x"857D797A", x"7C797677", x"6E6E6E6E", x"6C696A6C",
									 -- x"6D6D6D6E", x"6E6D6B6A", x"6F6C6B6C", x"6B68686B", x"6866676A", x"6E6D6B6A", x"6F707170", x"6E6C6661",
									 -- x"65686A69", x"66636465", x"68676A6C", x"6B6C6D6A", x"6B6B6966", x"676B6B68", x"6867696A", x"696B6D69",
									 -- x"6A68696A", x"696A6A66", x"676E726F", x"6C6D6F6E", x"75787876", x"787D7D7A", x"7C828480", x"80858581",
									 -- x"8581848D", x"8E89888E", x"908F8D8C", x"8E918F8C", x"8B898685", x"85878888", x"88888888", x"88888684",
									 -- x"82838485", x"85868788", x"86898A8A", x"8A8A8885", x"87868485", x"8987868A", x"8D8C8B8C", x"8E8E8C8A",
									 -- x"908F8E8D", x"8D8D8D8C", x"90959591", x"949B9D99", x"9B9B9A9B", x"9B9D9E9F", x"A0A0A0A0", x"A0A0A0A0",
									 -- x"A0A2A2A2", x"A2A4A5A5", x"A1A4A7A6", x"A3A2A6AA", x"A9A7A3A6", x"ADAAA8B0", x"ADABAAA9", x"ABADAFB0",
									 -- x"95989A9C", x"9C9D9FA0", x"A0A1A2A3", x"A3A4A5A6", x"A9A8A9AA", x"AAA9A9AA", x"A9A8A8AB", x"ACABAAAB",
									 -- x"B2B1B0B1", x"B2B4B3B2", x"B6B5B5B6", x"B8B9BABA", x"BCBCBDBE", x"BFBEBDBB", x"BEBEBEBD", x"BCBBBBBA",
									 -- x"BABBBBBB", x"BBBBBBBC", x"BFBEBEBF", x"BFBEBEBF", x"BDBDBEBE", x"BDBCBBBB", x"BCBBBAB8", x"B5B2AFAD",
									 -- x"A8A8A7A5", x"A4A4A6A7", x"A4A5A6A7", x"A8AAACAD", x"AEADADAF", x"B3B5B4B2", x"B2B0AFAF", x"B1B0AFAE",
									 -- x"AFAFAFAF", x"B0B0B0AF", x"ABABABAA", x"A7A4A2A1", x"A1A3A6A7", x"A7A6A6A6", x"A3A4A6A6", x"A7A9ABAC",
									 -- x"ABABABAB", x"ABAAA8A6", x"A8A7A6A5", x"A5A6A6A6", x"A2A2A3A3", x"A4A5A6A7", x"A6A5A5A5", x"A6A7A9AA",
									 -- x"AAAAA9A8", x"A7A7A8A9", x"A8A8A9A9", x"A9A9AAAB", x"ABAEAFAD", x"AEB1AFAC", x"ACACABAA", x"ABACABA9",
									 -- x"A7A6A6A5", x"A4A4A4A4", x"A3A4A5A6", x"A6A6A6A5", x"A9ABABAA", x"A9AAAAA9", x"A8A8A7A6", x"A8AAA9A7",
									 -- x"A6AAABA8", x"A8ACACA7", x"A9A9A9A8", x"A7A6A5A5", x"A5A4A3A2", x"A2A2A2A2", x"A2A0A0A0", x"A2A3A3A2",
									 -- x"A3A2A2A3", x"A3A2A2A4", x"A2A2A2A1", x"A0A1A4A7", x"A6A3A5AA", x"ABADAEAC", x"B0B0AFAF", x"AFB2B5B8",
									 -- x"BABDBFBF", x"BEC0C2C3", x"C5C4C3C4", x"C6C6C5C3", x"C4C5C5C3", x"C1C0C1C2", x"C1BEBDBD", x"BFC0BEBC",
									 -- x"BBBAB9B7", x"B6B3B1AF", x"AEAEAEAD", x"ADAEAEAE", x"ADADADAF", x"B0B1B0B0", x"ADADADAD", x"ADABA8A5",
									 -- x"A0A19F9A", x"97979591", x"91918F8E", x"8D8A8785", x"857F7876", x"797A7671", x"6F6E6F70", x"6D6A696B",
									 -- x"6C6C6B6C", x"6C6D6C6C", x"6E6A686A", x"6B69696A", x"6666686B", x"6C6B6A6A", x"6C6F706F", x"6E6B6763",
									 -- x"65696B6A", x"67656566", x"67666A6D", x"6C6D6D69", x"6E6D6964", x"65696865", x"67686B6A", x"66676A68",
									 -- x"6C696867", x"64666B6C", x"65686C6F", x"6F6F7072", x"78797875", x"777B7C7B", x"7C7F8282", x"807F8082",
									 -- x"84888987", x"898E8F8C", x"93928F8E", x"9092918D", x"8586898A", x"88868483", x"8A878584", x"84848281",
									 -- x"83828182", x"84858585", x"87888784", x"82838687", x"87868385", x"8A8A8687", x"8F8B8786", x"878A8C8E",
									 -- x"908E8C8B", x"8C8D8D8E", x"8D949591", x"91989C9A", x"98989797", x"999B9D9F", x"9F9FA0A0", x"A1A1A1A2",
									 -- x"A3A3A2A1", x"A4A7A7A5", x"A5A4A3A6", x"A9A9A6A3", x"A8A8A4A6", x"ACA9A9B3", x"ACABAAAA", x"ABACADAE",
									 -- x"93979B9D", x"9D9E9FA0", x"A2A3A4A5", x"A5A6A7A7", x"A8A7A8A9", x"A9A8A9AB", x"ADA9A7A9", x"AAAAABAD",
									 -- x"B0AFADAD", x"B0B3B2B0", x"B4B4B5B6", x"B8B9B9B9", x"BBBBBBBC", x"BEBEBDBC", x"BEBEBDBC", x"BBBBBABA",
									 -- x"BABBBBBB", x"BBBBBCBD", x"BEBDBCBD", x"BDBCBDBE", x"BEBFBFBE", x"BDBBBBBB", x"BCBBBAB9", x"B7B4B0AE",
									 -- x"AAA9A7A5", x"A3A2A2A2", x"A2A4A5A5", x"A4A5A9AD", x"AFAEABAB", x"ADB1B2B0", x"AEABAAAC", x"AFAFADAC",
									 -- x"ACACACAC", x"ADADADAC", x"AAAAA9A8", x"A5A3A1A1", x"9EA1A5A5", x"A4A3A3A5", x"A1A2A3A4", x"A5A6A9AB",
									 -- x"A8A8A8A8", x"A9A8A7A6", x"A6A6A5A4", x"A4A3A3A3", x"A2A3A3A3", x"A2A3A4A6", x"A4A3A4A7", x"A9A8A8A8",
									 -- x"A9A9A8A7", x"A6A7A8A9", x"A9A8A8A9", x"A9A8A9AB", x"ACADAEAE", x"AFB0AFAD", x"ADACAAAA", x"ABABAAA8",
									 -- x"A7A6A5A4", x"A4A3A3A3", x"A5A5A6A6", x"A6A5A4A3", x"A7A8A9A7", x"A7A8A9A8", x"A6A7A7A7", x"A8A9A9A7",
									 -- x"A8A9A9A8", x"AAADACA9", x"ABAAAAAA", x"AAA9A7A6", x"A6A5A4A4", x"A4A4A3A3", x"A3A1A0A1", x"A3A5A3A1",
									 -- x"A4A2A2A3", x"A4A3A3A4", x"A2A3A3A1", x"9F9FA2A5", x"A7A4A8AC", x"ACAEB0AF", x"B1B2B4B6", x"B6B7B8B8",
									 -- x"B8BCBFBF", x"BEC0C2C4", x"C4C3C2C5", x"C8C9C8C5", x"C4C5C5C4", x"C2C1C3C5", x"C4C2C0BF", x"C0C0BFBD",
									 -- x"C1BFBCBA", x"B7B3B2B2", x"B0B1B2B1", x"B0B0AFAE", x"B4B3B2B3", x"B5B5B4B2", x"B4B2AFAD", x"ADACABAA",
									 -- x"A5A4A09C", x"99989593", x"9392908E", x"8C898684", x"827E7775", x"797C7870", x"716F6E70", x"6E6A6869",
									 -- x"6A6A6A6B", x"6C6D6E6D", x"6A676669", x"6C6B6968", x"6465686A", x"69676768", x"6A6C6C6C", x"6C6D6C6A",
									 -- x"66676664", x"63646566", x"66636567", x"66686965", x"6C6B6865", x"65676765", x"69696A67", x"61636767",
									 -- x"6667696A", x"68666668", x"6B696A6D", x"6E6E7175", x"79787776", x"76787A7B", x"7E7E8285", x"837D7F85",
									 -- x"87868687", x"898C8F90", x"8E8F8F8F", x"90908D88", x"88888887", x"84828487", x"8C878483", x"85848382",
									 -- x"84828080", x"81828383", x"86888987", x"85858587", x"83878787", x"89878689", x"888A8B8A", x"86868A91",
									 -- x"918E8C8B", x"8C8C8E8F", x"8C939795", x"94989A98", x"97979797", x"999C9EA0", x"9D9E9FA0", x"A1A2A2A1",
									 -- x"A5A4A2A2", x"A6A9A9A7", x"A7A6A5A5", x"A6A6A5A5", x"A9A8A7A7", x"A9A7A8AF", x"A9AAABAC", x"ACADADAD",
									 -- x"9395989B", x"9D9F9F9F", x"A2A3A5A6", x"A6A7A7A8", x"A7A7A8A9", x"A9A8AAAC", x"ACA9A9AB", x"AAA8A9AC",
									 -- x"ACADADAD", x"AFB1B1AE", x"B1B2B3B5", x"B7B8B8B8", x"BABABABC", x"BEBFBEBC", x"BFBEBCBA", x"B9B9B9BA",
									 -- x"BABBBBBB", x"BABABCBD", x"BBB9B9BA", x"BABABBBD", x"BDBFBFBF", x"BDBCBBBC", x"BBBABAB8", x"B7B4B0AE",
									 -- x"AAA9A6A4", x"A3A2A1A0", x"9FA1A2A2", x"A1A2A7AA", x"AAABA9A7", x"A7A9ABAB", x"A8A7A7AA", x"ACABAAAA",
									 -- x"A8A8A8A8", x"A9A9A9A8", x"A7A7A6A4", x"A2A1A1A1", x"A0A1A2A2", x"A1A1A2A3", x"9FA1A2A2", x"A2A3A6A9",
									 -- x"A6A6A6A6", x"A6A6A5A4", x"A3A4A4A5", x"A4A3A2A1", x"A5A4A2A1", x"A1A1A1A1", x"A3A2A4A8", x"AAA9A8A8",
									 -- x"A8A8A8A8", x"A7A8A9AA", x"A9A8A8A9", x"A8A7A8AB", x"ACABACAE", x"B0AFAEAE", x"AEACABAB", x"ABABA9A8",
									 -- x"A6A5A5A4", x"A4A3A3A2", x"A5A5A6A6", x"A6A5A4A3", x"A5A7A8A7", x"A7A8A8A8", x"A6A8AAA9", x"A9A9A9A8",
									 -- x"A9A9AAAA", x"ABABACAC", x"ADAAA9A9", x"ABABA9A6", x"A6A5A5A6", x"A6A5A4A3", x"A4A3A3A3", x"A5A5A4A2",
									 -- x"A5A3A2A4", x"A5A3A3A3", x"A4A4A4A3", x"A2A1A3A4", x"A8A6AAAF", x"AEB0B3B3", x"B3B5B8BA", x"BABBBBBB",
									 -- x"B9BCBEBE", x"BFC1C2C2", x"C3C4C5C7", x"C9CACAC9", x"C6C6C5C5", x"C6C6C6C6", x"C7C5C3C1", x"C1C1C0BF",
									 -- x"C1BFBDBC", x"B9B5B4B5", x"B3B4B4B3", x"B2B2B1AF", x"B8B7B7B7", x"B8B8B8B8", x"B8B5B2AF", x"AFAEAEAD",
									 -- x"A8A5A2A0", x"9D999695", x"9493918F", x"8C8A8684", x"817C7878", x"7B7B7774", x"736E6C6D", x"6D6A6869",
									 -- x"69696A6B", x"6C6D6C6C", x"6A6A6967", x"68696866", x"63646667", x"67646465", x"68686768", x"6A6C6B67",
									 -- x"68686664", x"65686867", x"6A666768", x"686B6C69", x"69686869", x"68676667", x"68676866", x"62656967",
									 -- x"63696A6C", x"6F686164", x"6E6E6E6D", x"6C6E7072", x"79777779", x"7876787C", x"7F7F8287", x"85818286",
									 -- x"89818088", x"8B878990", x"8C8F9090", x"91908D8A", x"8C898683", x"8080858B", x"8A858285", x"87878584",
									 -- x"83838280", x"7E7F8284", x"8787898B", x"8B898684", x"81868886", x"87868589", x"84888D8E", x"8985888E",
									 -- x"8F8C8A8B", x"8C8B8D8F", x"8F929595", x"96979796", x"96969899", x"9B9C9D9E", x"9A9B9D9F", x"A0A09F9E",
									 -- x"A3A3A2A2", x"A4A7A8A7", x"A5A6A7A4", x"A1A1A5A9", x"AAA7A8A9", x"A8A8A9A8", x"A8AAACAD", x"ADADACAC",
									 -- x"93939598", x"9D9F9F9D", x"A1A3A4A5", x"A6A6A6A7", x"A7A7A9AA", x"AAAAABAE", x"A8A9ACB0", x"ADA7A6AA",
									 -- x"ACAFB0B0", x"B1B3B3B1", x"AFB0B2B4", x"B7B8B8B7", x"BAB9B9BB", x"BEBFBEBD", x"BFBEBBB9", x"B8B8B8B9",
									 -- x"B7B8B8B8", x"B7B7B9BB", x"BAB8B8B9", x"BABABBBD", x"BCBEC0C0", x"BEBDBCBC", x"BABAB9B8", x"B6B3B0AD",
									 -- x"A9A7A5A4", x"A4A3A1A0", x"9B9C9D9D", x"9D9FA3A5", x"A1A5A8A5", x"A3A3A5A6", x"A5A5A7A9", x"A9A7A7A9",
									 -- x"A5A5A5A5", x"A6A6A6A5", x"A4A4A3A1", x"A09FA0A0", x"A4A3A1A0", x"A0A0A0A1", x"9FA0A1A1", x"A0A1A4A7",
									 -- x"A7A6A5A5", x"A5A4A3A1", x"A1A3A5A6", x"A5A4A2A1", x"A3A09E9F", x"A1A3A3A2", x"A5A3A3A7", x"A9A9A9AA",
									 -- x"A7A8A8A8", x"A9A9AAAB", x"ABAAA9AA", x"AAA8AAAD", x"ACAAABAF", x"B0AEADAF", x"B0AEACAC", x"ACABAAA9",
									 -- x"A5A5A4A4", x"A4A3A3A3", x"A3A3A4A5", x"A5A5A4A4", x"A6A8AAA9", x"A9A9A8A7", x"A8ABADAC", x"AAAAAAA9",
									 -- x"A9AAABAC", x"ABA9AAAE", x"ADAAA7A7", x"A9ABA9A6", x"A4A4A5A6", x"A7A7A6A4", x"A4A5A6A6", x"A6A5A4A4",
									 -- x"A5A3A3A4", x"A5A3A2A2", x"A6A5A4A4", x"A5A5A5A4", x"A5A4A9AE", x"AEB0B4B5", x"B6B8B9BA", x"BBBCBDBF",
									 -- x"BEBFC0C0", x"C2C4C3C1", x"C7C8CACA", x"C9C8C7C7", x"C8C6C5C7", x"CACBC8C5", x"C7C6C4C3", x"C2C1C1C1",
									 -- x"BDBCBBBB", x"BAB6B6B7", x"B6B8B8B6", x"B5B6B5B3", x"B8B9BABA", x"BABABCBE", x"B7B6B4B3", x"B3B1AFAE",
									 -- x"ACA7A5A5", x"A39D9999", x"96949290", x"8D8B8886", x"847E7B7D", x"7C757274", x"746E696B", x"6C696869",
									 -- x"6A6A6B6C", x"6C6B6A68", x"6D6E6B65", x"62656666", x"63626365", x"65636262", x"66656466", x"696A655E",
									 -- x"62626161", x"63666460", x"67646568", x"696B6C69", x"6766686C", x"6B676668", x"66656768", x"676B6C68",
									 -- x"6C6E6765", x"6C686269", x"686E716D", x"6B6F7270", x"7977797D", x"7B76777D", x"7C7D8084", x"85838384",
									 -- x"86868685", x"878A8B89", x"898B8C8B", x"8B8C8B89", x"87868788", x"86838486", x"84807F83", x"87878482",
									 -- x"83858582", x"7E7E8388", x"89858283", x"86878583", x"82858484", x"87878687", x"87868686", x"8483878C",
									 -- x"8A888789", x"8B8B8B8E", x"90908F91", x"92949495", x"93949699", x"9A9A9A9A", x"999B9D9F", x"9F9F9E9D",
									 -- x"9EA0A1A0", x"A1A3A5A6", x"A6A29FA0", x"A3A6A7A6", x"AAA7A9AB", x"A9ABACA4", x"A9ABACAD", x"ADACABAB",
									 -- x"92969595", x"9B9F9F9F", x"9EA2A6A7", x"ABAEABA6", x"A9ABABA9", x"A8A9A9A8", x"A9AAAAAA", x"AAAAAAAA",
									 -- x"A8AAADB1", x"B3B2B1AF", x"B2B2B2B3", x"B4B6B7B7", x"B8B7B6B7", x"BABCBCBC", x"BBB9B8B6", x"B6B7B9BA",
									 -- x"B7B7B7B7", x"B7B7B7B7", x"B8B7B7B8", x"B9BBBBBC", x"B9BBBCBC", x"BCBCBBB8", x"B9B7B7BA", x"B9B5AFAB",
									 -- x"AAA7A3A0", x"A0A1A09E", x"9C9D9C99", x"989C9FA1", x"A8A3A1A4", x"A5A3A2A3", x"A2A2A1A1", x"A5A8A6A2",
									 -- x"A1A2A3A3", x"A3A3A3A3", x"A1A09F9F", x"9F9F9E9E", x"9FA0A1A2", x"A19E9D9F", x"A0A09F9E", x"9D9EA0A2",
									 -- x"A4A3A3A2", x"A2A2A2A2", x"A1A4A3A0", x"9FA1A2A0", x"9E9FA0A0", x"9F9FA0A1", x"A1A3A5A7", x"A7A7A8A8",
									 -- x"A9A8A7A6", x"A6A7A9AB", x"AEABAAAC", x"AEADABAA", x"A9AAABAD", x"AEAFAFAF", x"AFABA9AB", x"AEACA9A7",
									 -- x"A7A5A4A5", x"A5A2A1A2", x"A5A4A5A6", x"A6A4A5A7", x"A8AAA9A6", x"A5A9ACAB", x"AAABABAA", x"A9A9ABAC",
									 -- x"ABADAEAE", x"ADABABAB", x"AAABACAC", x"A9A8A8AA", x"A7A4A5A6", x"A3A5A7A5", x"A6A4A3A4", x"A6A7A6A5",
									 -- x"A8A5A2A2", x"A5A7A6A4", x"A4A4A1A0", x"A4A5A3A4", x"AAABACAE", x"B0B1B3B4", x"B7B8BABC", x"BDBEC0C2",
									 -- x"C5C5C5C5", x"C6C7C7C8", x"C8C7C8CB", x"CCCAC7C7", x"C8C7C6C5", x"C6C7C9CA", x"CAC7C4C3", x"C3C3C3C2",
									 -- x"BFBEBDBE", x"BEBCBAB7", x"BABDBEB9", x"B4B5B9BC", x"B8BCBEBC", x"BBBDBEBE", x"BFB9B8B7", x"B5B5B4AE",
									 -- x"AFADABA7", x"A29F9D9D", x"9A949092", x"928D8784", x"8383807B", x"77767471", x"726E6B6B", x"6B6B6B6B",
									 -- x"6A67676A", x"6C6A6868", x"63686A66", x"63646462", x"5E646562", x"6164635F", x"62656662", x"5F5F6161",
									 -- x"605E5D5E", x"61656869", x"63636968", x"696A6668", x"68666466", x"6A6D6C6A", x"67646A6D", x"68696A65",
									 -- x"6B696665", x"65666666", x"696D6F6F", x"6F727575", x"7E7B7878", x"78787A7C", x"85838085", x"8B84808A",
									 -- x"898A8681", x"858E8E87", x"878E8B89", x"888A8D87", x"88858384", x"85838384", x"867C8384", x"84868185",
									 -- x"86828081", x"7F7D7F83", x"85818282", x"7F838985", x"7D828484", x"84838790", x"8989888E", x"83858283",
									 -- x"89878588", x"8A8B8A89", x"8B8D8E90", x"93979897", x"9795969A", x"9C9A9999", x"98989A9D", x"9E9D9C9D",
									 -- x"9F9E9FA2", x"A4A3A3A4", x"A7A8A8A5", x"A1A1A4A9", x"A6A5A6A7", x"A4A2A6AC", x"ABAAA9A8", x"AAACABA8",
									 -- x"90949495", x"9CA0A1A2", x"A3A5A7A9", x"ABADADAC", x"ACADACAA", x"A8A9A9A8", x"A9A9A9A9", x"A8A7A7A6",
									 -- x"AAABADAF", x"B1B2B1B0", x"B0B1B1B2", x"B2B3B4B5", x"B7B7B6B6", x"B6B7B8B9", x"B9B8B6B5", x"B5B6B7B8",
									 -- x"B8B8B8B9", x"B9B8B8B8", x"B8B7B7B7", x"B9BABBBB", x"BBBCBDBB", x"BBBBBAB8", x"B9B8B7B8", x"B7B3AFAD",
									 -- x"A7A5A2A0", x"9F9E9C9B", x"9D9E9D9A", x"989A9C9C", x"A2A19F9D", x"9D9E9F9F", x"9E9E9D9C", x"9EA0A09D",
									 -- x"9F9FA0A0", x"9F9E9E9E", x"9F9E9E9F", x"A0A1A1A1", x"9F9F9FA0", x"9F9C9B9C", x"9D9D9C9C", x"9C9D9D9D",
									 -- x"9B9C9D9E", x"9FA1A1A2", x"A1A2A2A0", x"9FA0A09F", x"9F9F9E9F", x"A0A1A1A1", x"A2A4A6A7", x"A6A6A6A6",
									 -- x"ABAAAAA9", x"A9A9ABAC", x"ACABACAE", x"AEACABAB", x"ACACABAB", x"ABADAFB0", x"ADAAA9AB", x"ADABA8A7",
									 -- x"A9A6A5A6", x"A6A4A3A4", x"A3A2A3A5", x"A5A3A4A6", x"A9AAA9A7", x"A7AAACAC", x"ABABABAB", x"ABABACAD",
									 -- x"A8A9ABAB", x"AAAAAAAA", x"AAACADAB", x"A9A8A8A9", x"A5A3A6A7", x"A6A7AAA9", x"A7A6A4A5", x"A6A7A6A5",
									 -- x"A8A6A5A6", x"A8A8A7A5", x"A6A6A2A1", x"A5A6A6A9", x"AFB0B1B2", x"B4B6B9BB", x"B8BABCBD", x"BFC0C3C4",
									 -- x"C5C6C7C8", x"C8C9C9C9", x"CCCAC9C9", x"C8C7C8CB", x"C8C9CACB", x"CBCBCBCC", x"C8C6C4C3", x"C4C4C4C4",
									 -- x"C3C2C2C2", x"C1C0BFBE", x"BBBDBEBC", x"BBBBBCBB", x"BCBFC0BE", x"BDBFC0C1", x"C0BCBCBB", x"B6B5B4AF",
									 -- x"AEADABA8", x"A5A2A09F", x"A09B9593", x"928F8B89", x"8483807B", x"78777673", x"6F6C6A6B", x"6C6B6969",
									 -- x"6A676669", x"6A696868", x"64676763", x"62646564", x"63656460", x"5F636564", x"61656866", x"6362605E",
									 -- x"625E5B5D", x"63676764", x"64636968", x"68696668", x"69676565", x"67696969", x"6A696B69", x"656A6C64",
									 -- x"6E6D6B6B", x"6B6C6B6B", x"696A6C6F", x"6F6E7075", x"7C7F8282", x"7E7B7D81", x"87878180", x"8584848C",
									 -- x"8A898580", x"83898984", x"84898687", x"88898C88", x"87848488", x"8A888380", x"857D8283", x"81827E81",
									 -- x"82808083", x"817E7D80", x"83858989", x"86878986", x"82838181", x"8383848A", x"8785848A", x"83868383",
									 -- x"86858586", x"8A8D8D8B", x"8B8C8E90", x"94979794", x"96939294", x"97999B9D", x"9C9C9D9F", x"A09F9EA0",
									 -- x"9EA1A19E", x"A2A8A79F", x"A4A4A4A3", x"A3A4A7A9", x"A7A4A2A3", x"A5A5A5A5", x"AAABABAA", x"ABACABA9",
									 -- x"8E939394", x"9A9E9FA3", x"A6A7A9AB", x"ACACAEB1", x"AEAEADAB", x"AAABABAA", x"A9A9A8A8", x"A7A6A6A5",
									 -- x"ABABABAD", x"AFB0B1B1", x"AEAFB1B1", x"B1B2B3B5", x"B4B5B5B4", x"B3B3B5B8", x"B6B6B5B4", x"B4B5B5B6",
									 -- x"B6B7B8B9", x"B9B9B8B8", x"B8B7B6B6", x"B7B9BABA", x"BBBDBCBB", x"BABBBAB9", x"B9B8B6B6", x"B3AFACAC",
									 -- x"A5A4A3A2", x"A09D9B9A", x"9B9C9C9A", x"98999998", x"9C9F9D97", x"95999C9B", x"9B9C9B99", x"9A9B9B9A",
									 -- x"9D9D9D9C", x"9C9B9B9A", x"9C9B9C9D", x"9EA0A1A1", x"9F9D9C9C", x"9C999898", x"9998989A", x"9B9B9A98",
									 -- x"999A9B9D", x"9E9E9E9E", x"A09FA0A1", x"A09E9E9F", x"A09F9E9F", x"A1A2A2A1", x"A3A4A5A6", x"A6A5A5A5",
									 -- x"A8A9A9A9", x"A9A9AAAB", x"AAACAEB1", x"AFACABAB", x"AEADACAB", x"ABACADAE", x"ACABABAD", x"ADABA9A8",
									 -- x"AAA7A6A6", x"A6A5A5A6", x"A4A3A4A5", x"A6A5A6A8", x"AAA9A9A9", x"AAAAADB0", x"ADADADAD", x"AEAEADAD",
									 -- x"A9AAABAC", x"ACACACAD", x"ABACADAB", x"A9A8A8A8", x"A7A6A9AA", x"A6A7AAA9", x"A8A7A5A5", x"A6A7A6A5",
									 -- x"A5A6A6A7", x"A7A7A5A4", x"A6A7A4A2", x"A5A7A9AE", x"B1B2B2B4", x"B6B9BCBF", x"BCBDBFC0", x"C2C3C5C6",
									 -- x"C6C7C9CA", x"CBCBCBCB", x"CECECDCB", x"C8C7CACD", x"C7C8CACA", x"CBCBCBCC", x"C8C7C6C6", x"C6C6C5C4",
									 -- x"C4C4C4C3", x"C2C1C2C2", x"BFBFBEBE", x"C0C2C1BE", x"C1C3C3C2", x"C1C2C4C4", x"C1BFBFBD", x"B8B6B5B2",
									 -- x"AFAFAEAC", x"A9A5A3A1", x"A09E9994", x"918F8B88", x"84827F7B", x"79797774", x"6F6D6C6D", x"6E6C6A6A",
									 -- x"68666566", x"68676666", x"65656460", x"61646462", x"67656260", x"60616568", x"63656766", x"65635F5C",
									 -- x"5F5D5C5F", x"63666664", x"66646967", x"676A676B", x"6B686664", x"64656667", x"67696A66", x"656D7068",
									 -- x"6B6A6A6B", x"6C6C6B6A", x"6F6C6D72", x"716D6E74", x"767A7F81", x"7E7A7B7E", x"81858280", x"83848385",
									 -- x"8C898682", x"83868786", x"898B8689", x"8A878985", x"83838587", x"8784807E", x"807A8082", x"80828285",
									 -- x"7F7E8083", x"83818082", x"858B8D8B", x"8A888688", x"88868181", x"86868486", x"86838186", x"82848383",
									 -- x"82838384", x"898E8F8D", x"8C8D8E90", x"95989693", x"99969596", x"989B9EA1", x"9C9B9C9D", x"9E9E9FA1",
									 -- x"9EA2A29F", x"A1A7A6A0", x"A2A1A1A1", x"A3A6A7A8", x"A8A7A6A5", x"A7A8A6A2", x"A4A8ABAB", x"AAABABAB",
									 -- x"8E929292", x"96999BA1", x"A6A6A9AD", x"ACAAACB1", x"ADACABAB", x"ABACADAD", x"AAAAA9A9", x"A9A9A8A8",
									 -- x"AAA9AAAB", x"ADAFAFAF", x"ADAFB0B0", x"B0B1B4B6", x"B3B3B3B2", x"B2B2B5B6", x"B4B4B4B4", x"B4B4B4B4",
									 -- x"B3B4B6B7", x"B8B8B7B6", x"B7B6B5B5", x"B6B7B8B9", x"BABBBBBA", x"BABBBCBB", x"B9B8B6B4", x"B0ABA9A9",
									 -- x"A4A3A3A2", x"9F9C9B9B", x"989A9A98", x"98989897", x"9A9B9994", x"94969898", x"99999999", x"99999999",
									 -- x"99999899", x"99999998", x"9999999A", x"9B9C9D9D", x"9E9B9999", x"99979696", x"97969597", x"99999795",
									 -- x"98999A9C", x"9C9C9C9C", x"9E9D9EA1", x"A09C9B9E", x"9F9E9E9F", x"A0A1A2A2", x"A2A3A5A6", x"A6A6A6A7",
									 -- x"A5A6A7A8", x"A8A8A9AA", x"AAABAEB1", x"B1AEACAC", x"ACACADAD", x"ADACABAB", x"ACACACAC", x"ABA9A9A9",
									 -- x"A9A7A6A6", x"A6A5A4A4", x"A5A5A5A6", x"A6A6A7A9", x"A9A7A8AB", x"ACACAEB3", x"B0B0AFB0", x"B1B1AFAE",
									 -- x"ADAEAEAF", x"AFAEAEAE", x"ADADADAC", x"AAA9A8A8", x"A9A8AAAA", x"A6A6A9A9", x"A9A8A7A6", x"A7A7A7A6",
									 -- x"A5A6A7A7", x"A7A6A5A5", x"A6A8A6A4", x"A6A8ABB1", x"B0B1B3B5", x"B7BABDC0", x"C1C1C2C3", x"C4C5C6C6",
									 -- x"C8C9CBCC", x"CDCECECE", x"CECFD1D0", x"CECCCCCD", x"CBC9C7C7", x"C9CBCBCB", x"CACAC9C9", x"C8C7C6C5",
									 -- x"C4C5C5C3", x"C2C1C3C4", x"C5C3C0BF", x"C1C4C5C4", x"C4C6C7C6", x"C6C6C7C7", x"C3BFBFBD", x"B9B8B9B6",
									 -- x"B3B2B1AF", x"ACA7A3A0", x"9C9D9B95", x"918E8A85", x"84827F7C", x"7B797673", x"706E6D6E", x"6E6C6A6A",
									 -- x"66656464", x"65656464", x"64646260", x"6062615D", x"65636263", x"63616366", x"65656362", x"6262615F",
									 -- x"5B5E6161", x"61626669", x"67656967", x"676B6A6D", x"6B686565", x"65656666", x"66686866", x"686E6F6A",
									 -- x"67686869", x"6A6B6A6A", x"716D6C70", x"73727376", x"7A797A7D", x"7F7F7F80", x"80828383", x"83838282",
									 -- x"8A878584", x"8485878A", x"8C8B878C", x"8C878683", x"84858683", x"7E7C8084", x"7F7B7F82", x"82848687",
									 -- x"807F8083", x"84848689", x"8A8F8B86", x"86858489", x"8A878283", x"8A8A8686", x"87838385", x"81828383",
									 -- x"80828383", x"878E908D", x"908F8E8F", x"94989895", x"96969697", x"98999999", x"9A9A9A9B", x"9D9FA1A3",
									 -- x"9F9FA2A5", x"A39FA1A6", x"A2A3A2A2", x"A2A4A6A5", x"A8ABACA8", x"A5A6A6A5", x"A1A7ABAB", x"A8A7A8A9",
									 -- x"8F929090", x"949699A0", x"A3A5A9AE", x"ADAAABAF", x"ACABAAAB", x"ACADADAD", x"ABABABAA", x"AAAAAAAA",
									 -- x"A9A9AAAC", x"AEAFAEAE", x"AFAFAFAE", x"AEAFB2B4", x"B3B2B1B1", x"B2B3B4B4", x"B3B3B3B3", x"B3B3B3B3",
									 -- x"B1B2B4B6", x"B7B7B7B6", x"B6B5B3B3", x"B5B6B7B8", x"BABBBBBA", x"BABBBBBA", x"B9B8B7B5", x"B0AAA7A6",
									 -- x"A19F9E9E", x"9B98989A", x"97979795", x"95979897", x"9A959395", x"96959596", x"94959597", x"97969696",
									 -- x"95949495", x"96979796", x"97979798", x"999A9B9A", x"9C999797", x"97959494", x"96959394", x"97989795",
									 -- x"94959799", x"9A9B9B9B", x"9C9B9C9F", x"9E9A9A9C", x"9C9E9F9F", x"9E9EA1A3", x"A2A3A4A5", x"A6A6A6A7",
									 -- x"A5A6A8A9", x"AAABACAD", x"ABAAACB0", x"B2B1AEAC", x"ABACACAD", x"ADACABAB", x"ABABABA9", x"A8A8A8A9",
									 -- x"A8A8A8A7", x"A7A6A4A3", x"A4A5A5A4", x"A4A5A6A7", x"A9A7A9AD", x"AEADAFB3", x"B2B2B2B3", x"B5B5B3B1",
									 -- x"B1B1B0B0", x"AFAEADAC", x"AEAEAEAD", x"ABAAA9A9", x"A8A6A8A8", x"A5A7ACAC", x"A8A8A7A7", x"A8A8A8A8",
									 -- x"A8A9A9A9", x"A8A8A9AA", x"A7ABAAA9", x"ABABADB3", x"B2B4B7BA", x"BBBDBFC1", x"C4C4C5C6", x"C7C8C8C8",
									 -- x"CCCCCDCD", x"CECFD0D0", x"CFD0D1D1", x"D1D0CFCD", x"D1CCC8C9", x"CCCFCECC", x"CCCCCDCC", x"CBCAC8C7",
									 -- x"C8C8C8C6", x"C5C5C7C9", x"C9C6C4C3", x"C4C5C6C7", x"C6C7C9CB", x"CBCAC9C9", x"C7C1BEBC", x"BABBBBB7",
									 -- x"B6B5B3B1", x"ADA9A4A0", x"9C9E9D97", x"92908C87", x"8583817F", x"7D797572", x"716E6C6C", x"6B696869",
									 -- x"67666665", x"65656564", x"61606060", x"61615E5A", x"62606164", x"64606164", x"66636161", x"62636262",
									 -- x"5E606261", x"5F60656A", x"68656966", x"6669686B", x"6A666466", x"69686766", x"6969696B", x"6D6A6767",
									 -- x"6A6B6B6C", x"6D6D6E6E", x"6E6C6B6D", x"72787977", x"7B7A7A7B", x"7D7D7F80", x"86818082", x"80808388",
									 -- x"87848283", x"8383868A", x"8887848B", x"8D878684", x"8786847F", x"7D7F8488", x"83807F82", x"81818380",
									 -- x"81818284", x"8586888A", x"8C8F8882", x"8586868B", x"87868385", x"8A898586", x"87858786", x"82808485",
									 -- x"82848585", x"898E908E", x"928F8C8C", x"91969896", x"9697999A", x"9A9A9A9A", x"9C9C9C9D", x"9EA2A4A6",
									 -- x"A2A0A2A6", x"A4A0A1A6", x"A3A6A6A3", x"A1A3A5A5", x"A5A8A9A5", x"A3A5A6A5", x"A4A9ACAA", x"A6A4A4A4",
									 -- x"8F908F90", x"95979AA0", x"A1A4AAAD", x"ADABACAE", x"AEACABAC", x"ADACABAA", x"ACACABAA", x"A9A9A9A9",
									 -- x"A9A9ABAD", x"AFAFAEAE", x"B1B0AEAC", x"ACADAEAF", x"B4B2B0B0", x"B2B3B2B1", x"B2B2B3B3", x"B3B3B3B3",
									 -- x"B2B3B4B5", x"B6B6B6B6", x"B4B3B2B2", x"B3B5B7B8", x"B9BBBBBA", x"BABAB9B8", x"B9B7B6B4", x"B0AAA6A4",
									 -- x"A19E9B9B", x"99969698", x"96959492", x"92949593", x"96918F93", x"96939294", x"93929294", x"95959595",
									 -- x"94939393", x"95979796", x"95959596", x"989A9B9B", x"9A979695", x"95939293", x"95949293", x"94959695",
									 -- x"95969798", x"99999A9A", x"9A9A9B9D", x"9C9A999A", x"9A9C9E9D", x"9C9CA0A3", x"A2A3A4A5", x"A5A5A5A6",
									 -- x"A5A6A8A9", x"AAABADAE", x"ADAAAAAE", x"B1B1AFAE", x"ADACABAA", x"AAABACAD", x"ACADACAA", x"A9A9AAA9",
									 -- x"A8A9A9A9", x"A9A8A6A3", x"A5A6A6A4", x"A4A6A7A8", x"ABABACAE", x"AEAEAFB1", x"B3B4B5B6", x"B8B8B8B7",
									 -- x"B7B5B4B2", x"B1B0AEAD", x"B0AFAFAE", x"AEACACAB", x"ACA9A9A9", x"A6A8ABAA", x"A9A9A8A8", x"A8A8A9A9",
									 -- x"A9A9A9A8", x"A8A9ABAC", x"ABAFAFAF", x"B1B1B3B7", x"B5B8BCBE", x"BEBFC1C3", x"C7C7C7C9", x"CBCCCDCD",
									 -- x"CFCFCFCF", x"D0D1D2D2", x"D1D1D0CF", x"D0D2D1CF", x"D3CFCDCE", x"D2D3D0CC", x"CDCECFD0", x"CFCDCCCC",
									 -- x"CBCBCAC9", x"C8C9CBCD", x"CACACACB", x"CAC8C8C9", x"C9C9CCCE", x"CFCCCACA", x"CAC3BFBD", x"BBBCBBB7",
									 -- x"B7B5B3B0", x"AEAAA5A2", x"9F9E9A95", x"918F8D8A", x"87858482", x"7E797574", x"73706D6B", x"6967686A",
									 -- x"67686867", x"66676665", x"5E5E5E60", x"61615E5A", x"615F6061", x"615F6063", x"63616163", x"65646363",
									 -- x"65625E5E", x"60626464", x"66646764", x"63656366", x"68656569", x"6B696868", x"6869696D", x"6F6A666A",
									 -- x"6B6C6D6D", x"6D6D6E6F", x"73737170", x"73787874", x"787B7E7E", x"7A777A7F", x"817B7E83", x"807D8183",
									 -- x"85848283", x"8485878A", x"8A8A878C", x"8C868683", x"86827E7E", x"82868481", x"82817E81", x"7E7D827D",
									 -- x"82838485", x"85858586", x"8B8C8986", x"888B8B8D", x"88888788", x"8A888587", x"86848987", x"84808788",
									 -- x"8586878A", x"8D8F9090", x"928F8C8B", x"8F949694", x"95969797", x"989B9E9F", x"9F9F9F9E", x"A0A2A4A5",
									 -- x"A5A5A3A2", x"A5A9A6A0", x"A4A7A7A4", x"A2A4A7A7", x"A7A4A2A2", x"A6A9A8A5", x"A3A7A9A8", x"A7A6A6A6",
									 -- x"8D8E8E91", x"9798999E", x"A1A5A8A9", x"AAACAEAE", x"B0ADACAE", x"AEACA9A8", x"ABAAAAA9", x"A8A9A9AA",
									 -- x"A8A9AAAB", x"ADAEAEAD", x"B1AFADAD", x"AEAEADAC", x"B0B0B0B0", x"B0B0B0B0", x"B2B2B1B1", x"B2B2B2B2",
									 -- x"B3B3B4B4", x"B4B4B4B3", x"B3B2B0B1", x"B2B5B7B8", x"B7B9BBBB", x"BABAB8B6", x"B7B4B2B1", x"AEA9A5A3",
									 -- x"A29D999A", x"98959395", x"9292918F", x"90929290", x"92909091", x"92929293", x"94918F92", x"94959595",
									 -- x"94939191", x"93949392", x"93939395", x"97989999", x"98979595", x"93908F91", x"92929292", x"92939494",
									 -- x"97979797", x"98989898", x"989A9B9A", x"999A9998", x"999B9C9B", x"9B9C9FA2", x"A0A1A2A3", x"A3A4A5A6",
									 -- x"A5A6A7A8", x"A9AAABAC", x"AEACABAC", x"AEAEAEB0", x"ADACABAA", x"AAAAACAC", x"ABACACAB", x"AAABA9A7",
									 -- x"A7A8A9A8", x"A8A9A8A5", x"A5A7A7A5", x"A5A8AAAA", x"ABADAFAF", x"B0B1B2B2", x"B6B7B8B9", x"BABABABB",
									 -- x"BBBAB7B6", x"B5B4B2B0", x"B1B1B0B0", x"AFAFAEAD", x"B1ADACAC", x"AAABABA7", x"AAAAAAA9", x"A9A8A9A9",
									 -- x"A9A8A7A8", x"A9AAACAD", x"AFB2B2B2", x"B6B7B8BC", x"BABDC0C1", x"C1C1C4C6", x"CBCBCBCD", x"CFD1D2D1",
									 -- x"D1D1D2D2", x"D3D3D3D3", x"D2D4D3D1", x"D1D3D4D3", x"D3D1D0D1", x"D3D3D2D0", x"CFD1D2D2", x"D1D0CFCF",
									 -- x"CCCBCACA", x"CCCED0D1", x"CFCECDCF", x"CFCDCCCD", x"CDCCCED0", x"D0CDCBCB", x"CAC4C2C0", x"BDBCBCB8",
									 -- x"B8B5B2AF", x"ADAAA6A3", x"A09C9895", x"918D8B8A", x"87868482", x"7C767475", x"73706E6C", x"6A68686A",
									 -- x"66686967", x"66666664", x"605F5E5F", x"5F5F5E5E", x"5E5F6060", x"60606061", x"605F6063", x"64626162",
									 -- x"64615D5C", x"5F626363", x"62616562", x"61636063", x"6665686C", x"6B67686B", x"666C6B6B", x"6F6C6A6F",
									 -- x"6B6C6E6F", x"6E6D6D6D", x"76777878", x"76747475", x"7C7E8080", x"7C797C82", x"79788084", x"7F7E807C",
									 -- x"83838282", x"84888989", x"8C8D898B", x"89858784", x"82818182", x"85858079", x"7E828083", x"7E7C8583",
									 -- x"84848484", x"84848686", x"87888A89", x"888A8D8C", x"898A8788", x"8A888689", x"85828885", x"85818888",
									 -- x"8685878D", x"8F8F9093", x"9191908F", x"91939391", x"90929392", x"93969A9B", x"9D9FA09F", x"A0A2A4A3",
									 -- x"A7A8A7A6", x"A7A9A7A3", x"A7A9A7A4", x"A4A8A9A8", x"A9A5A3A6", x"AAAAA8A6", x"A3A4A5A5", x"A6A9A9A7",
									 -- x"8C8D8D92", x"9898979A", x"A1A4A6A5", x"A6ABAEAE", x"B1AEADAF", x"AFACA9A8", x"A9A9A8A8", x"A9AAABAC",
									 -- x"A7A7A8A9", x"ABACACAC", x"B0AEADAE", x"B1B1AFAC", x"ABADAFAF", x"AFAFB0B1", x"B1B1B1B0", x"B1B1B2B2",
									 -- x"B3B3B3B2", x"B2B1B1B1", x"B2B1B0B0", x"B2B4B7B8", x"B4B7BABB", x"BBBBB9B6", x"B4B0ADAC", x"ABA7A3A1",
									 -- x"A09A9697", x"96918F8F", x"8F8F8E8D", x"8F91908E", x"8E92928F", x"8F939493", x"95908C8E", x"91939394",
									 -- x"918F8D8C", x"8D8E8C8B", x"92929293", x"95969797", x"97969694", x"918D8D8F", x"90909191", x"91919293",
									 -- x"92929394", x"95979898", x"969A9B98", x"989A9997", x"9999999A", x"9A9C9EA0", x"9E9FA0A2", x"A3A4A5A6",
									 -- x"A6A7A8A8", x"A9AAABAC", x"AFADACAC", x"ABABAEB1", x"ABACACAC", x"ACABAAA9", x"A6A8A9A8", x"A8A8A6A2",
									 -- x"A5A7A7A6", x"A6A9A8A6", x"A3A5A5A3", x"A4A7A9A9", x"A9ADB0AF", x"B1B5B6B4", x"B9BBBCBB", x"BAB9BABB",
									 -- x"BCBAB8B7", x"B6B5B4B2", x"B2B1B1B1", x"B1B0AFAE", x"B0ACADAE", x"AEAFAEA9", x"ABABABAA", x"A9A8A8A9",
									 -- x"AAA9A9AA", x"ACADAEAF", x"B0B3B3B3", x"B8BABBBF", x"BFC1C4C4", x"C3C4C7CA", x"CFCFCFD0", x"D2D4D4D3",
									 -- x"D2D3D4D5", x"D5D5D4D3", x"D2D6D8D5", x"D3D4D5D5", x"D5D5D4D3", x"D2D3D5D7", x"D2D4D5D4", x"D2D1D0D0",
									 -- x"CECDCCCD", x"D0D3D4D4", x"D5D1CECF", x"D0D0D1D2", x"D1CFCFD1", x"D1CDCBCB", x"C7C4C4C3", x"BEBDBDBA",
									 -- x"B9B6B1AE", x"ACA9A5A3", x"A09B9898", x"958E8988", x"8684837F", x"79737376", x"706E6C6B", x"68676769",
									 -- x"64676765", x"64656462", x"64625F5E", x"5D5E5F60", x"5B5E6162", x"61615F5D", x"5F5D5D5F", x"605F6062",
									 -- x"5E5E5E5D", x"5D5F6366", x"5F5E6362", x"62646163", x"65676B6D", x"6964676D", x"69726F69", x"6C6C6B6F",
									 -- x"6E707374", x"73716F6F", x"6E70767B", x"7871737A", x"7B787676", x"77787A7D", x"7C7D8281", x"7B818680",
									 -- x"7F807F7F", x"83888987", x"888A8686", x"85848886", x"80868A89", x"85817D79", x"7F868688", x"807C8888",
									 -- x"86858381", x"8184888B", x"86858A89", x"83868C89", x"87878484", x"87868589", x"86828784", x"86818786",
									 -- x"8482858D", x"908E8F94", x"91939494", x"9494928F", x"96999A98", x"979A9B9B", x"9C9FA0A0", x"A1A4A5A4",
									 -- x"A8A7ABAE", x"A9A2A4AD", x"AAAAA7A3", x"A5AAABA7", x"A9A7A8AA", x"A9A5A4A6", x"A6A5A4A3", x"A4A6A5A2",
									 -- x"92909094", x"97999B9D", x"9F9FA0A2", x"A5A8ABAB", x"ADADADAD", x"ADACACAC", x"A8A7A7A7", x"A5A4A5A8",
									 -- x"A8AAAAAA", x"ACAEACA8", x"AAACADAC", x"ABADADAC", x"AFAFAFAE", x"ADADAFB0", x"B0B0B0B2", x"B2B0AFB0",
									 -- x"AEAEB0B3", x"B2B0B1B4", x"B0AEAEB1", x"B3B3B3B5", x"B7B8B9BA", x"BAB9B7B6", x"B1AFACAA", x"A8A6A2A0",
									 -- x"9C999997", x"9190908E", x"8F8F9090", x"8F8E8D8C", x"91908F8E", x"8F919292", x"8F8F8F90", x"91919090",
									 -- x"8F8D8A89", x"8A8B8B8B", x"8A8E908F", x"90939493", x"95969490", x"8F90908F", x"9190908F", x"90919292",
									 -- x"92909092", x"93939598", x"9B9C9C9B", x"9A999999", x"989A9C9C", x"9B9C9EA1", x"9D9FA1A2", x"A1A3A5A8",
									 -- x"A9A9A8A8", x"A9A9AAAA", x"ADAEAFAF", x"ADACACAD", x"AFAEACAB", x"ACABAAA9", x"A7A8A8AA", x"AAA9A6A3",
									 -- x"A7A8AAAA", x"AAA9A8A8", x"A8A8A6A4", x"A5A9AAA9", x"A9ADB1B3", x"B5B6B6B5", x"BABBBCBC", x"BDBFBEBB",
									 -- x"BDBDBAB8", x"B9BAB9B5", x"B6B5B3B2", x"B1B0B1B1", x"B1AFAEAE", x"AFAFAEAD", x"AAABACAB", x"AAA9A9AA",
									 -- x"ABACADAC", x"ABAAAAAA", x"ACB0B4B5", x"B7BABCBD", x"BDC0C4C5", x"C8CBCDCD", x"CCCFD2D3", x"D3D4D7D9",
									 -- x"D4D5D5D5", x"D5D6D7D7", x"D3D6D7D5", x"D4D7D8D6", x"D6D7D7D4", x"D4D5D6D6", x"D5D6D6D5", x"D6D8D7D4",
									 -- x"D1D0D0D2", x"D4D6D6D6", x"D8D7D5D5", x"D6D7D7D7", x"D3D4D4D5", x"D5D2CDC9", x"CAC6C2BF", x"BDBAB9BA",
									 -- x"B7B6B3AF", x"AEACA8A2", x"A09B9792", x"8F918E84", x"8487867E", x"78767673", x"726E6C6D", x"6E6C6B6B",
									 -- x"6E686567", x"68656465", x"61606164", x"625D5C5E", x"605C5C60", x"605D5C5F", x"5D5D6164", x"6262625E",
									 -- x"61605F5F", x"6162605D", x"64605F62", x"605C5F67", x"61656969", x"6A6B6A69", x"6E6D6E6E", x"6D6B6C6E",
									 -- x"7374726E", x"6C6F7172", x"71707476", x"767B7C72", x"7C797573", x"76797976", x"7D797D7C", x"827C8081",
									 -- x"8584817F", x"80838484", x"838E8D83", x"848F8D7F", x"84848584", x"83818181", x"81828388", x"8A858288",
									 -- x"8A878383", x"85878989", x"8B8B8988", x"8C92928F", x"9088858A", x"8D8A8687", x"898A8685", x"88848186",
									 -- x"8787888A", x"8D919496", x"96959697", x"97969697", x"9A9C9C99", x"989DA0A0", x"A39F9EA2", x"A9ABA8A6",
									 -- x"ACABABAB", x"ACACABA9", x"A9ACACA9", x"A9ADADAA", x"ABACACA8", x"A6ABACA4", x"A4A9A5A1", x"A6A8A5A5",
									 -- x"93929296", x"9999999A", x"9F9FA1A4", x"A7A9AAAA", x"ACACACAD", x"ACABABAA", x"A9A7A7A7", x"A7A6A7A8",
									 -- x"A9A8A7A6", x"A8ACADAC", x"AAACACAB", x"AAABABAB", x"ACACADAD", x"ADAEAFB0", x"AEACABAD", x"AFAFAFAF",
									 -- x"AFAEB0B1", x"B0AEAFB1", x"B1AEADAE", x"AFAFB0B2", x"B5B5B5B6", x"B8B8B6B3", x"B1AEABA8", x"A5A29E9C",
									 -- x"98959593", x"8F8F908E", x"8E8C8C8F", x"8E8C8C8D", x"8D8C8C8D", x"8E8F9090", x"8E8E8F90", x"9291908E",
									 -- x"8F8D8A89", x"89898989", x"898C8D8D", x"8E909090", x"94969490", x"8D8E8E8E", x"8F8F8F8F", x"8F8F8E8E",
									 -- x"8E8E8F91", x"92929599", x"97989999", x"99989898", x"989A9C9D", x"9D9D9FA0", x"A1A1A1A0", x"A0A2A6A9",
									 -- x"A9A9A9AA", x"AAABABAB", x"ADAEAFAF", x"AEAEADAD", x"ACABAAAA", x"AAAAA9A8", x"A9A9A8A9", x"A9A8A6A4",
									 -- x"A6A7A9A9", x"A9A8A7A7", x"A8A8A7A7", x"AAACACA9", x"ACAFB3B4", x"B6B9BAB9", x"BBBEBFBF", x"BEBEBEBD",
									 -- x"BEBEBDBA", x"BABCBAB8", x"B6B6B4B3", x"B3B3B4B5", x"B1B0AFAF", x"AFAFAEAD", x"ACADADAD", x"ABABABAC",
									 -- x"ABABABAB", x"ABABABAA", x"B2B5B7B7", x"B7BABCBD", x"C1C4C7C9", x"CBCECFCF", x"D1D3D5D7", x"D7D6D7D7",
									 -- x"D8D8D8D8", x"D7D6D6D6", x"D6D8D8D8", x"D7D9D9D9", x"D8D9D8D6", x"D5D6D7D6", x"D8D8D8D7", x"D7D9D8D5",
									 -- x"D5D5D5D7", x"DADBDBDA", x"DAD9D8D9", x"DADADAD9", x"D9D8D8D7", x"D7D4D0CD", x"CBC7C2BF", x"BDBABABA",
									 -- x"B6B6B4B0", x"ADABA6A1", x"A09C9893", x"90918F87", x"8185847D", x"79787876", x"74706D6E", x"6F6E6C6B",
									 -- x"6C666365", x"65636263", x"5E5E6064", x"64605F62", x"615D5C5E", x"5F5D5D61", x"5C5B5E60", x"5F61615F",
									 -- x"605F5E5D", x"5D5E6062", x"605F6164", x"63606063", x"65676866", x"65676969", x"6F6E6E6F", x"6D6B6C6E",
									 -- x"71747370", x"6D6F7375", x"73747575", x"767B7B76", x"73747676", x"78797775", x"7778787B", x"7B7C7C7F",
									 -- x"7E808383", x"83838586", x"81898B85", x"858A8983", x"81828383", x"8281807F", x"7D83827F", x"83878685",
									 -- x"86888C8D", x"8B87878B", x"93908E8E", x"8D8C8C8C", x"908C898B", x"8B888686", x"8D8B8786", x"88868486",
									 -- x"8B8A8A8C", x"91949695", x"9D9A9898", x"9797999B", x"9A9C9D9D", x"9D9EA0A0", x"A3A1A2A6", x"A9AAA9A8",
									 -- x"ACACACAC", x"ADADADAC", x"ABAEAEAB", x"ABADACA9", x"A8A8A9AA", x"AAAEAEA7", x"A8AAA8A5", x"A7A7A5A5",
									 -- x"93929498", x"9A9A9999", x"9D9EA1A4", x"A7A8A8A7", x"ABABACAC", x"ACAAA9A8", x"A8A6A6A7", x"A9A8A7A7",
									 -- x"A9A8A6A5", x"A7ABACAC", x"AAABABAA", x"A9ABABAB", x"AAABACAC", x"ACADAEAF", x"AEAAA8AB", x"AEAFAEAE",
									 -- x"AEAEAEAF", x"AEADADAE", x"B0AEACAC", x"ADADAEB0", x"B3B1B1B3", x"B6B7B4B1", x"B1AEAAA6", x"A3A09C99",
									 -- x"96939291", x"8D8D8F8E", x"8D8B8A8C", x"8C8A8A8C", x"8888898B", x"8C8D8D8D", x"8E8D8E90", x"91918E8B",
									 -- x"8E8C8988", x"87888888", x"898B8C8C", x"8C8E8F8E", x"8E90918E", x"8D8E9091", x"8E8F9091", x"91908E8D",
									 -- x"8D8D8F91", x"91929599", x"94959798", x"98989898", x"98999B9D", x"9E9F9F9F", x"A2A2A3A2", x"A2A3A6A8",
									 -- x"AAAAAAAB", x"ACACADAD", x"AEAEAEAF", x"B0B0AFAE", x"ADACACAC", x"ACACABAA", x"AAA9A8A7", x"A8A8A7A7",
									 -- x"A7A8A9AA", x"A9A8A8A8", x"AAAAABAC", x"AEB0AEAB", x"AFB2B5B6", x"B8BCBEBF", x"BEC1C4C2", x"C0C0C1C1",
									 -- x"C0C1C0BE", x"BDBDBDBC", x"B9B8B7B6", x"B6B6B7B7", x"B2B2B1B0", x"AEADADAE", x"AEAEAEAE", x"ADADADAD",
									 -- x"AEACABAB", x"ADAEAEAE", x"B4B7B8B8", x"B9BCBFC0", x"C4C8CBCC", x"CED1D2D2", x"D5D6D8D9", x"DAD9D7D5",
									 -- x"D9DADAD9", x"D8D7D6D6", x"D8D7D9DA", x"DAD9DADC", x"DADBDAD8", x"D7D8D8D7", x"DADADAD9", x"DADBDAD9",
									 -- x"D7D7D8DA", x"DCDDDDDC", x"DDDDDDDE", x"DEDEDDDC", x"DDDBD9D7", x"D6D4D1CF", x"CBC7C2C0", x"BDBBBABB",
									 -- x"B8B8B6B1", x"ACA7A29E", x"9E9C9B97", x"92928F88", x"8487857F", x"79787876", x"75706E6F", x"71706D6B",
									 -- x"6B666363", x"63616162", x"60606164", x"63605F61", x"615E5C5D", x"5D5C5E61", x"5B595B5E", x"5E60625F",
									 -- x"5F5F5F60", x"5E5D6167", x"5F616263", x"64646363", x"696B6B6A", x"6A6D7071", x"6F6F6F6F", x"6E6D6E71",
									 -- x"6F727371", x"6E6F7477", x"73777571", x"74767676", x"6E727677", x"78777573", x"7479777D", x"78807E81",
									 -- x"7B808586", x"84828488", x"8185898A", x"88878789", x"82848585", x"83807E7D", x"7E848380", x"84888684",
									 -- x"86888D92", x"908A898C", x"93909091", x"8F8B8C91", x"91908E8B", x"8A898888", x"8A898B8B", x"87868B8E",
									 -- x"8E8C8C8F", x"94979695", x"9F9C9A9A", x"9A9A9B9E", x"9C9DA0A4", x"A4A3A2A3", x"A5A6A9AB", x"ACABABAD",
									 -- x"AEAFAFAF", x"AFAEAFAF", x"AFB1B2AF", x"AEB0AFAC", x"ACA8A9AC", x"ACADACA7", x"A9A7A8A8", x"A5A4A5A4",
									 -- x"91929498", x"9A9B9B9B", x"9B9C9EA1", x"A4A6A6A5", x"AAABACAC", x"ABAAA8A7", x"A5A4A5A7", x"A7A6A5A6",
									 -- x"A9A9A8A8", x"A9AAA9A8", x"A8AAABA9", x"AAACADAD", x"AAABACAC", x"ACABACAC", x"ADABA9AB", x"ACACACAC",
									 -- x"ACACACAD", x"ADADADAE", x"ADACABAC", x"ADAEAFB0", x"B0AFAFB1", x"B3B4B3B1", x"B2AFABA7", x"A4A19D9B",
									 -- x"97939190", x"8C8C8E8C", x"8D8D8B89", x"88888887", x"8686888A", x"8C8C8B8B", x"8E8D8C8D", x"8F8F8D8A",
									 -- x"8B898887", x"87878889", x"88898A8B", x"8B8C8D8D", x"8A8C8E8D", x"8C8D9092", x"8E8F9091", x"91918F8F",
									 -- x"8E909292", x"91919498", x"94959697", x"98999A9A", x"9A9A9B9C", x"9E9F9F9E", x"A0A2A4A6", x"A6A6A6A7",
									 -- x"ACABABAB", x"ABACADAE", x"AFAEAEAF", x"B0B0AFAD", x"AEAEAEAE", x"AEAEADAC", x"A9A9A8A8", x"A9A9AAAA",
									 -- x"AAABACAC", x"ABABAAAA", x"ACADAFAF", x"B0B0B0B0", x"B2B5B7B7", x"BABEC1C2", x"C1C4C6C5", x"C4C4C5C4",
									 -- x"C2C3C2C1", x"BFBFBFBF", x"BEBDBBB9", x"B8B7B7B7", x"B3B4B3B1", x"AFADADAE", x"AEAEAEAE", x"AEADADAD",
									 -- x"AFADAAAB", x"AEB0B1B0", x"B2B6B8BA", x"BCC0C4C5", x"C6C9CCCE", x"D0D3D4D4", x"D8D7D8D9", x"DBDAD7D4",
									 -- x"D7D8D9D9", x"D8D7D7D7", x"D7D6D8DB", x"DBD9DADD", x"DCDDDDDA", x"D9D9DAD9", x"DADBDBDC", x"DDDEDEDE",
									 -- x"DADADADB", x"DCDEDEDE", x"E1E1E1E1", x"E1E0DFDE", x"DEDCD9D7", x"D5D3D0CE", x"CBC7C3C0", x"BEBCBCBD",
									 -- x"B8B8B6B2", x"ACA7A3A1", x"9E9D9D9A", x"93918E87", x"87888680", x"7B797877", x"74706E6F", x"71716E6B",
									 -- x"6B676464", x"63626163", x"62616162", x"625F5E5F", x"61605E5D", x"5C5C5E60", x"5C595B5D", x"5E60615E",
									 -- x"5C5D6064", x"635F6166", x"62636260", x"62666866", x"66686A6A", x"6A6B6D6E", x"6D6C6C6C", x"6C6B6E72",
									 -- x"6F717271", x"6F6F7275", x"72787570", x"73737276", x"73757675", x"76767472", x"7478787B", x"7A838281",
									 -- x"80828586", x"82808489", x"83868A8D", x"8B89898C", x"85868786", x"85838281", x"8385868A", x"8B878489",
									 -- x"8C87888F", x"918E8D8F", x"8F8F8F91", x"91909194", x"9192908C", x"8B8E8D8B", x"8C888B8D", x"888B8F8D",
									 -- x"8F8F8F91", x"95969695", x"9A999A9C", x"9D9C9C9E", x"9F9FA3A9", x"ABA8A7A9", x"AAABADAF", x"AFAEAFB2",
									 -- x"B1B2B3B3", x"B1B0B0B1", x"B1B3B3B1", x"B1B1B0AE", x"B0AAAAAD", x"AAAAABAB", x"AAA4A7AA", x"A4A1A4A4",
									 -- x"90929496", x"989A9B9C", x"9A9A9B9E", x"A1A4A5A6", x"A9AAABAC", x"ABAAA8A7", x"A3A4A7A8", x"A6A4A5A8",
									 -- x"AAAAAAAB", x"ABA9A7A6", x"A7A9AAA9", x"A9AAABAB", x"AAABACAC", x"ABABACAC", x"AAAAABAD", x"ACAAAAAC",
									 -- x"ACACACAB", x"ACADADAD", x"AAABABAC", x"ADAEAEAD", x"AEAFB0B0", x"B1B1B2B3", x"B3B0ACA8", x"A5A19D9B",
									 -- x"9792908F", x"8B8B8D8A", x"8B8E8D86", x"85898984", x"86878889", x"8B8B8A89", x"8D8C8A8B", x"8C8C8B89",
									 -- x"89898887", x"86878888", x"84858687", x"88888A8B", x"8C8D8E8D", x"8B8A8C8E", x"8F8F8F8F", x"8F8E8E8D",
									 -- x"8E909191", x"90919394", x"94959696", x"97989A9C", x"9D9C9B9B", x"9D9E9F9F", x"A0A2A5A7", x"A8A9A9A9",
									 -- x"AEADABAA", x"AAABADAF", x"B0AFAFAF", x"B0B0AFAD", x"ADADAEAD", x"ADACACAC", x"AAAAABAB", x"ABABACAC",
									 -- x"ADAEAFAE", x"AEADADAD", x"AEAFB0AF", x"ADADB0B4", x"B5B7B8B9", x"BBBFC2C3", x"C3C4C5C5", x"C6C8C7C5",
									 -- x"C5C5C4C3", x"C1C0C0C1", x"C0BFBEBC", x"BAB8B7B7", x"B6B6B5B2", x"AFAEAEAF", x"AFAFAFAF", x"AFAEAEAE",
									 -- x"ADAAA8A9", x"ACAFB0B0", x"B2B6B9BB", x"BEC2C4C5", x"C7CBCED0", x"D2D5D7D7", x"DBDAD9DA", x"DBDAD7D4",
									 -- x"D6D7D9D9", x"D9D8D8D8", x"D7D6D8DC", x"DCDADBDE", x"DDDFDEDC", x"DBDBDBDA", x"DCDCDDDE", x"DFDFE0E0",
									 -- x"DFDEDEDE", x"DFE0E2E3", x"E5E5E4E3", x"E2E1E0E0", x"E1DEDCD9", x"D7D5D1CF", x"CAC6C3C1", x"C0BEBDBE",
									 -- x"B7B6B4B1", x"ADAAA8A8", x"A19E9D99", x"928F8D89", x"8586847F", x"7C7B7B7A", x"75726F6F", x"70716E6B",
									 -- x"6B686664", x"63626263", x"5F5F5F60", x"60605F60", x"6162615F", x"5D5D5D5D", x"5D5A5C5E", x"5D5E5F5C",
									 -- x"595A5E62", x"63606062", x"64656360", x"62686A69", x"6A6A6B6A", x"68676869", x"6A696867", x"66676A6F",
									 -- x"71717171", x"71717172", x"70777572", x"76757378", x"75747474", x"76787673", x"75757774", x"7C7E807B",
									 -- x"807F8184", x"8482858B", x"8487898A", x"8B8B8A88", x"85868787", x"87878889", x"84888A8C", x"8C88878D",
									 -- x"908B8A8E", x"91909093", x"90939390", x"9094938E", x"9192908D", x"8E91908C", x"928A898C", x"8D919087",
									 -- x"90919495", x"96979798", x"9A999A9C", x"9D9D9E9F", x"A2A1A5AB", x"ADABABAD", x"AFAEAEB0", x"B1B1B3B5",
									 -- x"B3B4B5B5", x"B4B3B4B5", x"B3B4B3B2", x"B0B0AFAD", x"B0AAA9AB", x"A8A8ADB1", x"ACA6A8AB", x"A4A1A4A3",
									 -- x"91939494", x"95979999", x"9A9A9A9D", x"A0A3A6A7", x"A9A9AAAB", x"AAA9A8A7", x"A3A6A9AA", x"A6A3A5A9",
									 -- x"AAA9A8A9", x"A9A8A8AA", x"A7A9AAA8", x"A7A8A8A7", x"A9AAABAB", x"ABABACAD", x"AAABAEAF", x"ADABACAF",
									 -- x"ACACACAB", x"ACADACAA", x"AAABABAB", x"ACADACAA", x"ACAEAFAF", x"AFAFB1B3", x"B2B0ACA8", x"A4A09B98",
									 -- x"94908E8D", x"8B8C8D8A", x"898D8B85", x"84888884", x"87878888", x"898A8988", x"8C8B8988", x"88888888",
									 -- x"89898886", x"85858586", x"84848587", x"8788898C", x"8C8B8C8C", x"8C8B8C8D", x"9190908F", x"8E8D8D8C",
									 -- x"8C8D8E8E", x"8E909292", x"93939495", x"9697999B", x"9D9C9C9B", x"9C9E9FA1", x"A3A3A4A6", x"A8AAACAE",
									 -- x"B1AFADAB", x"ABADAFB0", x"B1B1B1B1", x"B1B0AFAE", x"AFAFAFAE", x"ADADADAE", x"AEAEAFAF", x"AEADADAD",
									 -- x"AFAFB0B0", x"AFAEAEAE", x"AEAFB0AF", x"ADACB1B6", x"B7B9BBBB", x"BDC0C2C3", x"C3C5C5C6", x"C8C9C8C6",
									 -- x"C8C7C5C5", x"C4C2C1C2", x"C0C0BEBD", x"BBBAB9B9", x"B8B7B5B3", x"B1B0B0B0", x"B1B0B0B0", x"B0B0AFAF",
									 -- x"ADABA9A9", x"ACAFB1B1", x"B4B8BCBD", x"BEC1C3C3", x"CACDD1D3", x"D5D8DADA", x"DFDDDCDC", x"DCDBD8D5",
									 -- x"D8D9DADA", x"D9D8D7D7", x"D6D7D9DC", x"DDDDDDDF", x"DDDFDFDD", x"DCDCDCDB", x"DEDEDFE0", x"E0DEDFE0",
									 -- x"E1E1E1E1", x"E1E2E4E6", x"E7E7E6E4", x"E2E1E1E1", x"E0DEDBD9", x"D7D4D0CE", x"CAC7C4C3", x"C1BFBDBE",
									 -- x"BBB8B4B1", x"ADAAA8A9", x"A59F9C96", x"908E8F8D", x"88878480", x"7C7A7A7A", x"78767370", x"70706E6B",
									 -- x"6A696766", x"64636363", x"62616060", x"60605F5F", x"60636360", x"5E5E5E5D", x"5D5B5D5E", x"5B5B5C5A",
									 -- x"5C5C5D5F", x"60616261", x"61646564", x"65686968", x"6C6B6A69", x"6867696B", x"6B696867", x"6666696D",
									 -- x"73717072", x"73727170", x"6D717374", x"75757476", x"71717274", x"787B7874", x"77747772", x"7B787C77",
									 -- x"7B797D85", x"8784858A", x"83868686", x"888B8983", x"8A8A8988", x"87878889", x"818C8C85", x"868C8E8E",
									 -- x"90929494", x"928F9194", x"91969590", x"9196948D", x"9292908F", x"9092908B", x"8A8B8E8E", x"8C8E9291",
									 -- x"93959899", x"999A9B9D", x"A09E9D9D", x"9E9FA1A4", x"A5A4A6A9", x"ACADAEAF", x"B2B0B0B2", x"B4B5B5B6",
									 -- x"B4B5B6B7", x"B6B6B7B7", x"B7B7B6B4", x"B2B1B0AF", x"B1ABAAAA", x"A6A6ACAF", x"ABA7A7A6", x"A2A0A1A0",
									 -- x"90929492", x"92949695", x"99999A9C", x"9FA2A4A5", x"A8A8A9A9", x"A9A9A8A8", x"A5A6A8A9", x"A6A4A5A8",
									 -- x"A8A6A6A7", x"A6A6A7AA", x"A7AAABA9", x"A8A8A8A6", x"AAAAABAA", x"AAAAABAC", x"ACACADAD", x"ACAAABAD",
									 -- x"AAABABAA", x"ABADACA9", x"ABACACAB", x"ABACACA9", x"ACACADAD", x"ADAEAFB1", x"AFADAAA7", x"A4A09A97",
									 -- x"948F8E8E", x"8C8D8E8B", x"8B8A8887", x"86848484", x"87878686", x"87888888", x"89898988", x"86858686",
									 -- x"87878785", x"84838485", x"86858688", x"8887898C", x"8B89898C", x"8D8D8D8E", x"908F8F8E", x"8E8D8D8D",
									 -- x"8B8C8C8C", x"8E91918F", x"90929495", x"9798999A", x"9B9C9C9C", x"9C9EA0A2", x"A4A4A4A6", x"A9ACAEAF",
									 -- x"B2B1B0AF", x"AFB0B1B2", x"B1B2B3B3", x"B2B1B1B1", x"B3B3B3B1", x"AFAFB0B2", x"B1B2B2B1", x"B0AFAFB0",
									 -- x"B0B1B1B1", x"B0AFAFB0", x"B0AFB0B2", x"B2B2B4B7", x"B9BBBEBE", x"C0C3C4C4", x"C5C7C9C9", x"C9CACAC9",
									 -- x"CCC9C6C7", x"C6C4C2C2", x"C0C0BFBE", x"BDBCBBBB", x"BAB8B6B4", x"B3B2B1B1", x"B1B0AFAF", x"B0B0AFAE",
									 -- x"ADACABAB", x"ACAFB2B3", x"B5B9BCBD", x"BEC2C4C5", x"CCCFD3D4", x"D6DADBDB", x"DEDEDEDE", x"DEDCD9D6",
									 -- x"D9D9D9D8", x"D7D6D6D6", x"D5D8DBDC", x"DDDFE0DF", x"DDDFDFDD", x"DCDDDDDC", x"DFDEDFE1", x"E0DEDEE0",
									 -- x"E1E2E3E3", x"E3E3E4E5", x"E5E6E7E6", x"E4E2E2E2", x"DEDCD9D6", x"D4D2CECC", x"CAC8C5C4", x"C2BFBCBC",
									 -- x"BEBAB5B2", x"AEAAA7A6", x"A39D9B98", x"9392928F", x"8E8C8883", x"7F7B7A7A", x"79797672", x"71717170",
									 -- x"6C6B6A69", x"67656564", x"66646261", x"6161605F", x"5F636460", x"5E60605E", x"5F5D5F5E", x"59595C5B",
									 -- x"5D5F5F5D", x"5E626361", x"5F626566", x"66666767", x"64646465", x"64636568", x"68686969", x"6968696C",
									 -- x"6E6E6F71", x"72707071", x"6E6E7174", x"73737472", x"70717273", x"76787673", x"75747576", x"77767779",
									 -- x"79777C85", x"86818187", x"85858687", x"898B8985", x"8E8E8D8B", x"89878787", x"858D8B83", x"878F918F",
									 -- x"92969996", x"93929393", x"90949693", x"93969592", x"91929393", x"9493908E", x"868E918D", x"8B8D939A",
									 -- x"9697999B", x"9C9E9FA0", x"A4A1A0A1", x"A2A3A5A8", x"A8A9A9AA", x"ACAFB0AF", x"B4B3B4B7", x"B9B9B9BA",
									 -- x"B8B8B7B8", x"B8B8B7B7", x"B8B7B5B4", x"B3B2B2B2", x"B0ABA9A9", x"A7A9AAA8", x"A6A7A39F", x"A0A09F9F",
									 -- x"8E919392", x"92939494", x"9898999B", x"9EA0A2A2", x"A7A7A7A8", x"A8A8A8A8", x"A5A5A6A7", x"A5A3A4A5",
									 -- x"A6A4A5A6", x"A6A4A5A7", x"A7AAACAB", x"ABABAAA8", x"ACACABAA", x"A9A9A9AA", x"ACA9A8A8", x"A8A6A6A7",
									 -- x"A7A9A9A9", x"ABAEADAA", x"ACADADAB", x"ABAEAEAC", x"ACABAAAA", x"ACADAEAE", x"ADABA9A7", x"A4A19C98",
									 -- x"95919090", x"8E8F8F8B", x"8E888689", x"87807F84", x"87858484", x"85878888", x"86888988", x"86848485",
									 -- x"84858584", x"83838486", x"86848486", x"8685878A", x"8E8B8A8C", x"8E8D8B8B", x"8A8B8B8C", x"8C8D8D8D",
									 -- x"8C8D8C8C", x"8F92918E", x"8F919497", x"99999A9A", x"989B9D9D", x"9D9EA1A3", x"A3A4A6A8", x"ABADAEAD",
									 -- x"B2B2B2B3", x"B3B3B4B4", x"B1B3B4B4", x"B3B2B3B4", x"B6B5B4B2", x"B0B0B1B3", x"B2B3B3B2", x"B1B1B2B3",
									 -- x"B2B2B3B2", x"B1B1B1B1", x"B1B0B1B5", x"B9B8B8B8", x"B9BDBFC1", x"C2C5C6C6", x"C7CBCECC", x"CBCBCCCC",
									 -- x"CECAC7C8", x"C8C5C3C2", x"C1C1C0BF", x"BEBDBCBB", x"BBB9B6B4", x"B4B3B3B2", x"B0AFAEAE", x"AFAFAEAD",
									 -- x"ACACABAB", x"ABADB0B3", x"B4B7BABC", x"BFC4C8CA", x"CDD0D3D4", x"D6D9DBDA", x"DBDCDEDF", x"DFDDDAD7",
									 -- x"D7D7D7D6", x"D5D5D5D6", x"D4D8DBDB", x"DCE0E0DE", x"DCDEDFDD", x"DDDDDDDC", x"DDDDDEE0", x"E0DEDFE1",
									 -- x"E1E3E5E6", x"E6E5E5E5", x"E4E5E7E7", x"E6E4E2E2", x"DEDCD8D5", x"D3D1CECC", x"CBC9C7C6", x"C3BFBCBB",
									 -- x"BBB6B2B2", x"B0ACA9A8", x"9D9A9B9D", x"9996938D", x"8F8D8986", x"82807F7F", x"797A7874", x"72747575",
									 -- x"6D6E6D6B", x"69686766", x"64636262", x"64656564", x"5F646460", x"5E616260", x"615F615F", x"59595D5E",
									 -- x"595E605C", x"5C60615D", x"60616466", x"65646668", x"6566686A", x"69656364", x"62636669", x"6968696B",
									 -- x"696A6D70", x"706E6E71", x"736F7477", x"73737470", x"73747371", x"70727271", x"6F717178", x"7275747C",
									 -- x"7B797C83", x"827C7D84", x"8886878A", x"8C8C8B8B", x"8C8D8E8E", x"8C8B8B8B", x"8B8B898A", x"90918F90",
									 -- x"95979693", x"94979691", x"91949797", x"95939496", x"90929698", x"97949293", x"93938B87", x"90949292",
									 -- x"9797989B", x"9EA0A1A1", x"A2A1A2A5", x"A7A7A8AA", x"ABADADAB", x"ADB2B2AF", x"B5B6B9BD", x"BDBCBCBD",
									 -- x"BCBAB9B9", x"B9B8B6B4", x"B3B2B1B0", x"B0B1B2B3", x"ABA7A6A8", x"AAAEADA6", x"A3A7A19C", x"A2A4A1A3",
									 -- x"8B909190", x"90949696", x"9998989B", x"9D9E9E9F", x"A3A5A6A5", x"A3A3A4A6", x"A4A5A5A4", x"A3A4A7AA",
									 -- x"A5A7A7A6", x"A6A6A6A4", x"A5A6A8A8", x"A9A9A9AA", x"ACAAA9A8", x"A9A9AAAA", x"A5A8ABAA", x"A7A6A8AB",
									 -- x"AAA7A7A9", x"ABAAAAAB", x"A7A9AAAB", x"ABABABAA", x"ABACACAA", x"A9AAACAD", x"ACA8A5A6", x"A5A09B99",
									 -- x"9894908D", x"8D8D8C8B", x"89888786", x"84838282", x"7F828585", x"84838384", x"87868785", x"82858783",
									 -- x"84828183", x"84838384", x"81838586", x"86858585", x"87888889", x"89898988", x"8A8C8D8C", x"8A898B8D",
									 -- x"8C8E8F8E", x"8D8D8E8F", x"8D8F9294", x"95969899", x"9C9D9D9E", x"9FA0A1A2", x"A1A2A5A9", x"ABACAFB3",
									 -- x"B5B7B8B7", x"B7B6B4B2", x"B5B6B5B3", x"B3B4B3B1", x"B6B5B4B5", x"B6B5B3B1", x"B2B2B3B4", x"B5B5B4B3",
									 -- x"B2B3B2B2", x"B1B2B3B3", x"B2B3B4B5", x"B6B8BBBC", x"BBBCBFC2", x"C2C2C6CA", x"CBCCCDCE", x"CDCDCCCC",
									 -- x"CECCC9C6", x"C6C7C6C4", x"C2C3C1BE", x"BEBFBEBB", x"BBBAB8B7", x"B6B5B3B2", x"AEAFAFAE", x"AEAFADA9",
									 -- x"A9A9AAAC", x"ADAEAFAF", x"B3B8B9BA", x"BEC0C3CA", x"CDD0D3D5", x"D6D7D8D9", x"DDDDDDDD", x"DDDBD9D6",
									 -- x"D6D7D7D5", x"D5D8D9D8", x"D8DADCDD", x"DDDDDEDE", x"DCDEE0DF", x"DDDCDEE0", x"DFE0E0DE", x"DEE0E1E0",
									 -- x"E1E3E4E5", x"E4E4E5E6", x"E7E8E8E8", x"E7E5E2E0", x"DFDEDBD6", x"D1CECDCD", x"CCC7C3C3", x"C3C0BDBC",
									 -- x"BBB7B3B2", x"AFAAA6A5", x"A29E9D9E", x"9C959294", x"908D8A86", x"817C7C7F", x"7E7B7774", x"73737272",
									 -- x"6D6D6A69", x"6A676568", x"65626164", x"64626264", x"65636260", x"605F5F5F", x"605C5A5D", x"5D5B5D61",
									 -- x"5C5C5B5C", x"5C5D5D5C", x"625E6066", x"66626165", x"61616264", x"64636260", x"66626367", x"66676A6B",
									 -- x"6667686A", x"6E706D68", x"6F737571", x"70727473", x"6D6A7073", x"7174766E", x"6D727273", x"76757476",
									 -- x"7A7C7F82", x"83848484", x"83868185", x"878E8989", x"8C8C8F92", x"918E8C8C", x"918E8D90", x"93949494",
									 -- x"98959599", x"9C9B9997", x"97999896", x"97959293", x"95939496", x"95919093", x"938E908F", x"9296969C",
									 -- x"9A98999E", x"A3A3A2A1", x"A1A8AAA7", x"A7ABADAB", x"B8B2B1B6", x"B9B6B7BA", x"B7B8BABC", x"BDBDBBBA",
									 -- x"BCBCBCBC", x"BCBAB7B4", x"B7B4AFAE", x"AEB0B0B0", x"AEA8A7A9", x"A9ABABA6", x"A3A4A5A5", x"A3A19E9C",
									 -- x"888C8F90", x"91939494", x"979A9C9A", x"9A9D9F9E", x"A0A2A3A3", x"A2A3A5A7", x"A6A6A6A5", x"A4A5A8AA",
									 -- x"A8AAA9A6", x"A4A5A6A7", x"A6A6A7A8", x"A8A8A8A8", x"AAA9A8A8", x"A9AAABAB", x"A6A9ACAC", x"AAA9AAAC",
									 -- x"A9A7A7A8", x"AAA9A9AA", x"A8A9AAAB", x"ABAAA9A8", x"A7A8A8A8", x"A7A7A8A9", x"AAA6A4A4", x"A29E9997",
									 -- x"95928F8D", x"8C8C8B89", x"89888887", x"86858484", x"81838484", x"83828283", x"84838584", x"8182837F",
									 -- x"82818285", x"85838283", x"83848585", x"85858585", x"86868787", x"87878686", x"898A8A8A", x"89898A8B",
									 -- x"8B8D8E8F", x"8E8E8F90", x"8F909293", x"94959798", x"9B9C9E9F", x"A0A1A3A4", x"A3A4A7AB", x"ADAEB1B5",
									 -- x"B7B9BCBC", x"BBBBB8B5", x"B8B8B6B4", x"B3B5B4B3", x"B6B5B4B4", x"B4B5B5B5", x"B3B4B5B6", x"B7B7B6B6",
									 -- x"B6B6B5B4", x"B4B4B6B7", x"B4B5B6B7", x"B8B9BABB", x"BEBDBFC2", x"C4C4C6C9", x"CBCCCECE", x"CECDCDCD",
									 -- x"CFCECBC9", x"C8C9C8C6", x"C1C2C2C0", x"C0C1C0BD", x"BCBBBAB9", x"B8B6B4B3", x"B1B1B0AE", x"AEAEADAB",
									 -- x"ACABAAAB", x"ACAEB1B3", x"B3B8BABB", x"BFC1C3C9", x"CCCFD2D4", x"D6D7D8D9", x"DBDDDEDD", x"DBD9D8D7",
									 -- x"D7D7D6D6", x"D6D6D6D6", x"D7D8DBDC", x"DDDDDEDE", x"DDDFE0E0", x"DFDEDFE0", x"E0E1E0DE", x"DEE0E0DF",
									 -- x"E1E3E5E6", x"E5E4E4E4", x"E6E5E5E5", x"E4E2E0DE", x"DEDDDAD5", x"D0CDCCCC", x"C8C7C4C0", x"BFC0BDB9",
									 -- x"B7B4B1B0", x"ADA9A5A4", x"A4A3A09D", x"9A979491", x"908D8B89", x"84807F80", x"7C7B7876", x"75757676",
									 -- x"70706D6B", x"6D6A686C", x"65686760", x"60656560", x"6463615F", x"5E5D5E5E", x"605D5C5E", x"5E5C5D60",
									 -- x"5959595A", x"5C5F6061", x"5E5F6263", x"62616162", x"60606060", x"60605F5E", x"63616569", x"65646565",
									 -- x"64666868", x"6A6B6B69", x"6C6D6E6E", x"6D6D6F71", x"6C6C716F", x"686D7676", x"70727172", x"76767476",
									 -- x"7A7C7E81", x"84868788", x"888D8A8C", x"8889858A", x"8A8A8B8E", x"8E909398", x"8F8D8D90", x"94959697",
									 -- x"9B979495", x"98999899", x"97979594", x"97979698", x"95939396", x"95919194", x"918F9699", x"9C9E9A9D",
									 -- x"999DA1A2", x"A1A0A2A5", x"A7ABACAA", x"AAAEB1B2", x"B7B6B6B9", x"B9B6B6B8", x"BDBDBDBE", x"BFBFBFBF",
									 -- x"BEBDBCBD", x"BEBDB9B6", x"B8B5B2B1", x"B3B4B4B3", x"ADAAABAD", x"ACABA8A2", x"A1A1A1A0", x"9F9F9F9F",
									 -- x"87888A8E", x"90919294", x"969C9E99", x"989D9F9E", x"A0A1A2A2", x"A2A3A5A7", x"A6A6A6A6", x"A5A5A7A9",
									 -- x"A6A9AAA7", x"A3A4A6A8", x"A7A6A6A7", x"A8A9A8A6", x"AAAAA9A9", x"AAAAA9A9", x"A8A9ABAC", x"ACABABAB",
									 -- x"A8A7A6A7", x"A8A8A8A9", x"AAAAAAAA", x"A9A8A7A6", x"A4A5A5A5", x"A4A4A4A5", x"A7A4A2A1", x"9F9B9795",
									 -- x"94928F8D", x"8C8B8987", x"87868686", x"85858585", x"82848484", x"82828283", x"81808282", x"7F7F7F7A",
									 -- x"80818385", x"84828182", x"82838383", x"82838485", x"84848585", x"85858484", x"87878787", x"87888888",
									 -- x"898B8D8E", x"8E8E9091", x"90919293", x"94969899", x"9D9E9FA0", x"A1A2A4A5", x"A5A7AAAE", x"B0B2B5B8",
									 -- x"B8BBBDBE", x"BDBDBAB7", x"B9B8B6B3", x"B3B5B5B4", x"B5B4B3B2", x"B2B2B4B6", x"B4B6B8B8", x"B8B8B9BA",
									 -- x"BAB9B8B6", x"B6B7B9BA", x"B6B7B8BA", x"BABABBBB", x"C1BFBFC2", x"C5C6C7C8", x"CBCCCECF", x"CFCECECF",
									 -- x"CFCECCC9", x"C9CAC9C6", x"C3C4C4C3", x"C3C3C1BF", x"BEBDBCBA", x"B9B7B5B4", x"B4B4B3B0", x"AEAEAFAE",
									 -- x"ADADACAC", x"ADB0B3B4", x"B4B9BCBE", x"C2C3C4C8", x"CBCED1D3", x"D5D6D7D8", x"D9DBDCDB", x"D8D6D6D7",
									 -- x"D8D5D5D7", x"D7D5D5D7", x"D8D9DBDD", x"DDDEDEDE", x"DFDFE0E0", x"E0E0E0E0", x"E1E1E1DF", x"DEDFE0DF",
									 -- x"DDDFE1E3", x"E3E2E1E0", x"E5E4E3E2", x"E1E0DFDE", x"DFDDDAD5", x"D0CDCBCB", x"C5C8C6BF", x"BCBFBDB7",
									 -- x"B4B1AFAE", x"ACA9A6A4", x"A2A3A09A", x"9A9C9A94", x"8F8C8988", x"8582807F", x"7B7A7876", x"75757677",
									 -- x"71706D6B", x"6C6A696D", x"676A6861", x"5F646460", x"6464625F", x"5D5C5D5F", x"5C59595B", x"5B58585A",
									 -- x"5B5A595A", x"5C5E5F60", x"5B606361", x"5F606160", x"6160605F", x"5E5E5E5E", x"61616667", x"62606161",
									 -- x"62666968", x"67686A6A", x"6866676B", x"6B696B70", x"6C6A6D6E", x"6D717572", x"74757272", x"76777577",
									 -- x"7B7C7D7F", x"80838587", x"888A888E", x"8989868B", x"8D8C8C8C", x"8D8E9398", x"92909093", x"96969596",
									 -- x"9F9B9797", x"99999A9A", x"999A9796", x"9A9B999B", x"97959597", x"96939497", x"93929A9C", x"9FA19DA0",
									 -- x"9DA3A7A5", x"A3A5A9AA", x"A8AAACAC", x"ADAEB2B5", x"B7BABDBD", x"BBB9B9B9", x"BFBFBFC0", x"C0C0BFBF",
									 -- x"C0BEBDBE", x"C0BFBCB8", x"B9B7B5B5", x"B6B6B5B3", x"ADABAEAF", x"ACA9A7A1", x"A3A2A09E", x"9E9FA1A2",
									 -- x"8986868A", x"8E8F9297", x"979B9C9A", x"999D9F9F", x"A3A3A3A3", x"A3A4A5A7", x"A5A5A6A5", x"A4A5A6A7",
									 -- x"A2A6A9A7", x"A5A5A6A6", x"A8A6A5A6", x"A9AAA8A7", x"A9A9A9A9", x"AAAAAAA9", x"A9A9A9AA", x"ABABAAA9",
									 -- x"A8A7A7A7", x"A8A8A8A8", x"AAAAAAAA", x"A9A8A6A5", x"A5A4A3A4", x"A3A2A3A4", x"A2A19F9E", x"9C999695",
									 -- x"95949290", x"8E8B8886", x"86868686", x"86868686", x"83848584", x"84838383", x"807F8181", x"7E7E7D7A",
									 -- x"7F818484", x"82808182", x"7E7F8080", x"80808283", x"82838384", x"84848383", x"85858485", x"86878787",
									 -- x"88898A8B", x"8B8C8F91", x"90919394", x"96999B9D", x"A1A1A2A2", x"A3A4A5A6", x"A8AAACAF", x"B1B4B8BB",
									 -- x"BABCBEBE", x"BEBDBAB7", x"B7B7B5B3", x"B4B6B6B5", x"B5B6B6B5", x"B3B2B3B4", x"B4B6B9B9", x"B8B8BABC",
									 -- x"BAB9B9B8", x"B7B7B9BA", x"B7B8BABB", x"BBBCBDBF", x"C1C1C1C3", x"C5C7C8C9", x"CBCCCECF", x"D0D0D0D1",
									 -- x"D0CFCDCB", x"CBCBCAC7", x"C6C6C6C5", x"C4C3C1BF", x"BFBEBDBB", x"BAB8B6B5", x"B5B6B5B2", x"B0B0B1B2",
									 -- x"ADADAEB0", x"B1B2B3B3", x"B5BABEC0", x"C4C5C5C9", x"CBCDD0D2", x"D4D5D6D6", x"D7D9DAD9", x"D7D6D6D8",
									 -- x"D7D4D4D9", x"D9D6D6DA", x"DBDCDDDE", x"DEDDDDDD", x"E0DFDFE0", x"E1E2E1E0", x"E2E2E1DF", x"DEDFDFDE",
									 -- x"DADBDEDF", x"E0E1E1E1", x"E4E3E2E1", x"E1E0DFDE", x"DEDDDAD6", x"D2CECBC9", x"C6C8C7C0", x"BCBCBBB7",
									 -- x"B4B2AFAE", x"ADAAA8A6", x"A3A39F9B", x"9C9E9C96", x"908C8886", x"8583817F", x"7E7D7C79", x"76747575",
									 -- x"71716D6B", x"6C6B6A6D", x"68666566", x"64616063", x"64646360", x"5E5D5F61", x"5F5D5C5D", x"5C5B5B5C",
									 -- x"5C5B5A5A", x"5C5D5D5D", x"5C5E6060", x"5F606060", x"6060605F", x"5E5D5C5D", x"62606263", x"5F5F6261",
									 -- x"61666968", x"6768696A", x"65646669", x"6A696B6F", x"6B6A6B6E", x"7174746F", x"76767372", x"7677777A",
									 -- x"7F7F7E7D", x"7D7F8285", x"8B85828C", x"8B8D8A8C", x"8F8F8F90", x"90909090", x"95949497", x"99989898",
									 -- x"A2A09F9F", x"9F9E9C9B", x"9B9E9C9B", x"9D9B999B", x"9B999999", x"9897979A", x"9B989B99", x"9AA0A1A7",
									 -- x"A2A4A3A2", x"A7AEAFAA", x"A6A7ACB0", x"B1AFB0B4", x"B9BDC0BF", x"BFC0BFBD", x"BDBFC2C3", x"C3C1BFBD",
									 -- x"C1C0BFBF", x"BFBFBEBD", x"BCB9B6B5", x"B5B5B2B0", x"AFADAEAD", x"A8A7A8A6", x"A7A4A09E", x"9D9D9EA0",
									 -- x"8785868A", x"8D8F9398", x"9A98989C", x"9E9E9FA2", x"A4A4A4A4", x"A4A4A5A6", x"A5A5A6A5", x"A5A5A5A6",
									 -- x"A4A6A7A6", x"A6A7A6A5", x"A8A6A5A7", x"A9ABAAA9", x"A6A6A7A9", x"AAACACAC", x"ABAAA9A8", x"A9AAA9A9",
									 -- x"A9A8A8A7", x"A8A9A9A8", x"AAA9A9A9", x"A9A8A7A5", x"A6A3A2A2", x"A1A0A1A3", x"9D9D9D9B", x"99989695",
									 -- x"94939290", x"8E8B8987", x"88888887", x"87868686", x"83848484", x"83828180", x"817E7F80", x"7D7D7E7C",
									 -- x"7F818281", x"7F7F8082", x"7D7E7F7F", x"7E7E7E7F", x"7F808182", x"82828282", x"84838384", x"85878787",
									 -- x"87888888", x"888A8D90", x"91929495", x"979A9D9E", x"A3A4A4A5", x"A5A6A8A9", x"ABADAEAF", x"B1B5BABD",
									 -- x"BEC0C0BF", x"BEBDBCB9", x"B8B8B7B6", x"B6B7B6B4", x"B5B7B9B9", x"B7B5B4B4", x"B3B6B8B8", x"B8B8BABC",
									 -- x"B9BABABA", x"B9B9B9B9", x"BBBBBBBB", x"BBBDBFC1", x"BFC2C4C4", x"C5C7C9CB", x"CACCCED0", x"D1D2D2D3",
									 -- x"D3D3D1CF", x"CFCFCDCA", x"CAC8C6C5", x"C4C3C2C1", x"C0BFBEBC", x"BBB9B7B6", x"B4B4B5B4", x"B2B1B1B3",
									 -- x"AFAFB0B1", x"B2B3B3B4", x"B6BCBFC2", x"C7C7C7CA", x"CCCDCFD2", x"D3D4D4D4", x"D8D8D7D8", x"D8D8D8D8",
									 -- x"D7D3D4D8", x"D9D5D6D9", x"DADBDDDE", x"DDDDDDDD", x"E0DFDEDF", x"E1E2E1DF", x"E2E2E1DF", x"DEDFDFDD",
									 -- x"DCDDDDDF", x"E0E1E2E2", x"E2E1E1E1", x"E1E0DEDC", x"D9D9D8D6", x"D3CFCBC9", x"C7C7C5C2", x"BDB8B7B8",
									 -- x"B5B3B1AF", x"AEACA9A6", x"ACA7A2A0", x"9F9D9A97", x"94908B87", x"86868482", x"8382807D", x"7A787777",
									 -- x"7475716E", x"6F6E6D70", x"6867686A", x"68626062", x"63636260", x"5E5E6061", x"5F5D5B5B", x"5A5A5B5C",
									 -- x"5959595A", x"5C5D5E5D", x"5E5A5A5F", x"615E5D5F", x"5D5E5E5E", x"5C5B5A5A", x"605E5F60", x"60636562",
									 -- x"62656768", x"68696967", x"66686967", x"676A6B6A", x"686D6F6C", x"6C6E7277", x"71757473", x"7576797E",
									 -- x"8282817F", x"7F808487", x"9189868F", x"8B8F8E8F", x"8E8F9093", x"96969492", x"9595979B", x"9D9E9FA0",
									 -- x"A2A3A3A3", x"A2A19F9D", x"9A9F9E9D", x"9C9A999D", x"9E9D9C9C", x"9B999A9B", x"A29E9F9A", x"9BA1A3A9",
									 -- x"A4A4A2A1", x"A8B1B1AB", x"AAAAAFB4", x"B5B3B4B8", x"BDC0C0BF", x"C1C4C4C0", x"C0C2C5C6", x"C6C4C2C2",
									 -- x"C2C2C1C0", x"BEBEBFC0", x"BDBAB7B5", x"B4B3B1AF", x"B0ADADAB", x"A6A6A8A6", x"A7A29F9D", x"9C9A9A9B",
									 -- x"8385898D", x"8F909396", x"9C97989F", x"A19F9FA3", x"A2A2A3A3", x"A4A5A5A6", x"A6A6A7A7", x"A7A6A6A6",
									 -- x"AAAAA7A4", x"A4A6A7A6", x"A8A7A6A7", x"A9ABABAA", x"A9A9A8A9", x"A9AAA9A9", x"ABAAA9A9", x"A9AAAAAA",
									 -- x"A9AAA9A8", x"A8AAA9A8", x"A8A7A6A7", x"A8A8A7A5", x"A5A19FA0", x"9F9D9D9F", x"999B9B99", x"97969696",
									 -- x"8F8F8F8E", x"8D8B8988", x"87868686", x"85858484", x"84848382", x"817F7E7D", x"827E7E7F", x"7C7C7E7D",
									 -- x"7F807F7D", x"7C7D7F80", x"7E7E7F7E", x"7D7C7C7B", x"7C7C7E7F", x"80808080", x"82828384", x"85868788",
									 -- x"87888887", x"87898C8F", x"92939597", x"989A9C9E", x"A3A4A6A7", x"A9AAACAE", x"AEB0B1B1", x"B3B8BCBF",
									 -- x"BFC0C0BE", x"BDBCBBB9", x"BBBCBBB9", x"B8B8B7B4", x"B3B5B7B8", x"B7B6B5B4", x"B4B5B7B7", x"B7B8BABB",
									 -- x"BBBCBDBC", x"BCBBBBBB", x"BFBEBDBC", x"BCBDBFC1", x"BFC3C5C5", x"C5C7CACC", x"CACCCFD1", x"D2D3D4D5",
									 -- x"D5D5D3D1", x"D1D0CDCA", x"CBC8C6C6", x"C5C3C3C3", x"C1C0BFBD", x"BCBBB9B8", x"B4B3B4B5", x"B4B2B1B2",
									 -- x"B4B3B2B1", x"B1B3B5B7", x"B8BDBFC2", x"C8C9C9CD", x"CDCECFD1", x"D3D4D3D2", x"D5D5D4D5", x"D6D7D6D5",
									 -- x"D7D4D4D7", x"D7D5D5D7", x"D7D9DBDC", x"DDDDDDDE", x"DFDFDEDF", x"E1E1E1DF", x"E2E2E1DF", x"DEDFDFDD",
									 -- x"DEDEDDDD", x"DEE0E0E0", x"DFDFDFDF", x"DFDEDCDB", x"D4D4D4D4", x"D3D0CDCA", x"C8C5C3C2", x"BEB8B7B9",
									 -- x"B5B4B2AF", x"AEADAAA7", x"ADA9A4A3", x"A19E9B9A", x"96938D88", x"86868583", x"8483807E", x"7D7B7978",
									 -- x"77787470", x"71716F71", x"686E6F69", x"6667645F", x"61605F5F", x"5E5F5F5F", x"5B5A5857", x"56575859",
									 -- x"5A5A595A", x"5A5B5B5A", x"5E57565C", x"5F5B5A5D", x"5C5D5E5E", x"5C5B5B5C", x"5E5C5E61", x"62666661",
									 -- x"63646566", x"68696866", x"696C6B67", x"666A6966", x"676D6E6D", x"70717073", x"6E737473", x"75777A81",
									 -- x"7F808181", x"8184888B", x"908B8B92", x"888E9294", x"92929394", x"989B9A98", x"9A9A9B9E", x"A0A0A1A3",
									 -- x"A2A3A3A1", x"A0A0A1A1", x"9DA1A09F", x"9F9FA0A5", x"9F9F9F9E", x"9D9C9D9E", x"A0A0A5A3", x"A2A5A2A5",
									 -- x"A9ABABA9", x"ABB0B2B1", x"B0B0B2B5", x"B6B6BABF", x"C1C2C1C0", x"C2C5C4C1", x"C5C6C6C5", x"C4C4C5C6",
									 -- x"C3C3C2C1", x"BFBEBFC1", x"BDBAB7B5", x"B5B4B2B0", x"AFACADAC", x"A7A5A5A3", x"A5A19E9F", x"9F9C9A9B",
									 -- x"81878C8E", x"8E919495", x"9B9A9CA0", x"A2A0A1A3", x"A1A2A3A4", x"A6A6A6A6", x"A6A6A7A7", x"A7A7A6A5",
									 -- x"ABABA8A4", x"A3A4A6A7", x"A7A7A7A7", x"A8A9AAAA", x"ACABAAA9", x"A8A8A7A7", x"A8A9AAAA", x"ABAAAAAA",
									 -- x"A9AAA9A8", x"A8AAA9A7", x"A7A5A4A5", x"A6A7A6A4", x"A39F9EA0", x"9F9B999A", x"96999A97", x"94949594",
									 -- x"8E8E8E8D", x"8B898887", x"86868585", x"85848484", x"86848281", x"80808080", x"807C7C7D", x"7A797B7A",
									 -- x"7D7D7C79", x"797B7C7C", x"7D7D7D7C", x"7B7A7B7B", x"7B7C7D7E", x"7F7F7F7F", x"80818384", x"84858788",
									 -- x"87888989", x"898A8D8F", x"9495989A", x"9B9D9FA0", x"A5A6A8A9", x"ABADAFB1", x"B1B4B5B5", x"B7BBBEC0",
									 -- x"BEC0C0BE", x"BDBDBBB9", x"BDBDBBB9", x"B8B9B9B7", x"B6B5B5B5", x"B6B6B5B5", x"B6B6B7B7", x"B8B9BABA",
									 -- x"BDBEBEBE", x"BDBCBCBD", x"C0BFBFBD", x"BDBDBFC0", x"C1C4C5C4", x"C5C8CACA", x"CACCCFD1", x"D3D4D5D6",
									 -- x"D6D6D4D2", x"D1D0CDC9", x"CDCAC8C8", x"C7C4C2C2", x"C2C1C0BF", x"BEBDBBBA", x"B7B5B5B6", x"B6B4B3B3",
									 -- x"B7B6B4B3", x"B3B5B6B8", x"B9BDBFC2", x"C9CBCCCF", x"CDCDCFD1", x"D3D4D3D2", x"D3D4D4D4", x"D4D4D4D4",
									 -- x"D7D6D6D6", x"D6D6D7D8", x"D7D9DBDD", x"DDDEDEDF", x"DFDFDFE0", x"E1E1E1E0", x"E2E2E1DF", x"DEDFDFDE",
									 -- x"DDDCDCDC", x"DDDEDEDD", x"DFDEDDDD", x"DDDDDCDB", x"D6D5D4D4", x"D3D1CECC", x"C7C7C5C2", x"BFBDBCBB",
									 -- x"B5B5B3B0", x"AFAFACA8", x"A8A8A5A1", x"9F9F9E9A", x"96948F8A", x"87888785", x"83817E7D", x"7E7D7A77",
									 -- x"77797571", x"71716F6F", x"6B706F67", x"63666662", x"62605F5F", x"60605F5D", x"5D5D5C5A", x"5A5B5B5C",
									 -- x"5D5B5958", x"57585858", x"5C59585A", x"5B5A595A", x"5B5D5E5D", x"5C5B5D5E", x"5F5E6061", x"61656662",
									 -- x"65666565", x"66696968", x"6C6B6A69", x"69696968", x"696E6D6F", x"7877706E", x"72767676", x"78797A7F",
									 -- x"7E818385", x"85878A8D", x"8D898B91", x"868E9493", x"94969796", x"96999B9B", x"A09FA0A1", x"A1A0A1A3",
									 -- x"A2A4A4A1", x"A0A2A4A5", x"A3A6A5A5", x"A8A7A5A6", x"A0A1A2A2", x"A1A1A2A2", x"9FA2ABAA", x"A9ABA6A6",
									 -- x"AEB0B1B0", x"AFB0B3B6", x"B3B5B6B7", x"B8BABEC1", x"C3C4C4C4", x"C4C5C4C4", x"C6C6C6C5", x"C3C2C4C6",
									 -- x"C5C4C2C2", x"C2C2C0BE", x"BCBAB7B7", x"B7B5B2B0", x"ADAAABAB", x"A7A6A5A1", x"A4A09EA1", x"A19E9C9D",
									 -- x"81888D8B", x"8B909597", x"999EA1A1", x"A0A1A2A3", x"A3A3A5A6", x"A8A8A7A6", x"A5A5A6A6", x"A7A6A5A3",
									 -- x"A6A8A9A6", x"A3A3A5A6", x"A7A7A8A7", x"A7A7A8AA", x"A9A8A7A7", x"A8AAABAB", x"A4A7A9AB", x"ABAAAAAA",
									 -- x"A9AAA9A7", x"A8A9A9A7", x"A6A4A3A4", x"A5A6A5A3", x"A29E9EA0", x"A09A9797", x"95989995", x"92929393",
									 -- x"8F8F8F8D", x"8A888685", x"88888888", x"88888787", x"87848280", x"80828485", x"7F7A7A7C", x"78767877",
									 -- x"7B7B7977", x"777A7A79", x"7A7A7979", x"78797B7D", x"7C7D7E7E", x"7F7F7F7F", x"7F818383", x"83848689",
									 -- x"87888A8B", x"8C8C8E90", x"95979A9C", x"9FA1A3A4", x"A7A8AAAB", x"ACAEB0B1", x"B2B6B9B9", x"BABDC0C0",
									 -- x"BFC1C2C1", x"C1C0BEBB", x"BBBBB9B7", x"B8BABAB9", x"BDBAB7B6", x"B6B8B8B8", x"B8B7B7B8", x"B9BABBBA",
									 -- x"BFBFBEBD", x"BDBCBDBE", x"BEBFBFBE", x"BEBFC0C1", x"C3C4C4C4", x"C6C9C9C8", x"CACCCFD2", x"D3D5D6D7",
									 -- x"D8D8D7D5", x"D3D2CECA", x"CFCCCBCB", x"C9C4C1C0", x"C2C1C0C0", x"BFBEBDBB", x"BCB9B7B8", x"B9B7B5B6",
									 -- x"B7B7B7B7", x"B7B7B6B6", x"BABEBFC2", x"C9CCCDD1", x"CCCDCED1", x"D4D5D4D3", x"D5D7D9D8", x"D6D4D5D6",
									 -- x"D7D8D8D6", x"D7DADBDB", x"DADBDDDE", x"DFDFDFDF", x"DFDFE0E0", x"E1E1E1E1", x"E1E2E1DF", x"DEDFDFDE",
									 -- x"DCDCDCDE", x"E0E0DFDE", x"E0DFDDDC", x"DCDCDCDC", x"DAD9D6D5", x"D3D1CECC", x"C7CAC8C2", x"C0C3C2BD",
									 -- x"B6B6B4B1", x"B0B1AEAA", x"A6AAA79E", x"9A9D9B94", x"9797938E", x"8B8B8A88", x"85817F7F", x"80807C79",
									 -- x"787B7772", x"73726F6F", x"6E6B6866", x"63616368", x"63615F60", x"61625F5C", x"5B5B5B5A", x"5A5A5A5A",
									 -- x"5B595655", x"56585B5C", x"5B5C5C5A", x"595A5A58", x"595A5B5A", x"59595C5E", x"6261615F", x"5D626664",
									 -- x"68686765", x"66696B6C", x"6D69696C", x"6C6A6A6C", x"6C747370", x"73737379", x"797C7A79", x"7C7B797C",
									 -- x"8285898A", x"89898B8E", x"928B8A90", x"8892938B", x"91969997", x"95989B9D", x"A09FA0A2", x"A2A2A4A6",
									 -- x"A2A5A7A5", x"A4A6A7A7", x"A5A8A8AB", x"AFABA39F", x"A2A4A5A5", x"A5A6A6A6", x"A4A7AFAD", x"ADB0ADAE",
									 -- x"B1AFAFB1", x"B1B1B2B5", x"B5B8BCBC", x"BDBFC1C2", x"C4C5C7C8", x"C7C6C6C8", x"C5C7C8C7", x"C5C3C3C4",
									 -- x"C7C4C2C3", x"C6C5C0BB", x"BBB9B8B8", x"B7B5B1AE", x"ACA8A8A8", x"A5A6A7A4", x"A29E9DA0", x"A19D9B9C",
									 -- x"82868A8D", x"8F909294", x"959AA0A2", x"A2A3A2A1", x"A4A4A4A5", x"A6A6A5A4", x"A7A5A4A5", x"A8A8A7A6",
									 -- x"A9A8A8AA", x"AAA7A6A8", x"A8A8A8A8", x"A7A7A9AB", x"AAA9A8A8", x"A8A9AAAA", x"A7ABAEAD", x"ADADADAC",
									 -- x"AAABA9A7", x"A6A7A7A6", x"A6A5A5A4", x"A4A4A3A2", x"A1A09E9E", x"9E9B9793", x"95949393", x"93939291",
									 -- x"908E8C8C", x"89868587", x"88878889", x"89888583", x"80838584", x"84848381", x"807C7878", x"77757678",
									 -- x"77777879", x"78787878", x"78777778", x"7877797B", x"7B7C7A7C", x"82827E7E", x"82838483", x"84868888",
									 -- x"8C8B8B8D", x"8D8E9195", x"95989B9D", x"9EA0A2A4", x"A8A8AAAC", x"ACADAFB3", x"B4B6B9BA", x"BBBDBFC1",
									 -- x"C2C3C3C1", x"C0C0BFBD", x"B9B9BABA", x"BABABABA", x"BBBAB9B8", x"B7B7B6B6", x"B9B8B8B9", x"BABCBBBB",
									 -- x"BDBDBDBC", x"BBBABCBE", x"BDBFC0C1", x"C0C1C2C3", x"C6C3C3C5", x"C5C5C7CA", x"CACCCFD1", x"D3D5D6D8",
									 -- x"D3D6D6D3", x"D1D2CFCB", x"CACAC9C8", x"C6C4C4C4", x"C3C1C0C0", x"BFBCBBBB", x"BBBABBBD", x"BCB9B7B8",
									 -- x"BAB9B8B7", x"B8B8B8B8", x"B9C1C5C6", x"C8CACBD0", x"CECECFD0", x"D2D4D4D4", x"D7D8D9D9", x"D9D9D9D9",
									 -- x"D7D7D8D8", x"D8DADBDD", x"DADCDEDF", x"DEDEDEDF", x"E0DFDEDF", x"DFE0DFDF", x"E1E2E1DF", x"DFE1E2E1",
									 -- x"DEDEDDDD", x"DEE0DFDC", x"DBDCDEDF", x"E0DEDBD9", x"DCD7D5D7", x"D4CDCDD1", x"CECAC7C7", x"C5C1BEBD",
									 -- x"B9B7B5B5", x"B6B5B2AF", x"AAA6A5A6", x"A29E9B96", x"9795928E", x"8F8F8B85", x"82818181", x"81818180",
									 -- x"79787674", x"71707070", x"6F6A6665", x"67686765", x"5F625D5E", x"5C595E5D", x"58595C5F", x"5E5A5859",
									 -- x"5B57575C", x"5C585658", x"595B5B58", x"56575959", x"5C5C5859", x"5E5B5960", x"61605F5F", x"61646667",
									 -- x"63696669", x"6964686B", x"6A6E6E6B", x"6A6D6E6C", x"6D6D6F75", x"79767882", x"7B7F807F", x"7F7D7C7F",
									 -- x"81868583", x"888D8D8E", x"93929293", x"95979694", x"94989997", x"999D9D9B", x"A1A1A1A2", x"A3A6A9AB",
									 -- x"AAABACAB", x"A9A8A9AB", x"AAAEB0AC", x"ACAEADA8", x"A7AAABA9", x"A7A8A9A9", x"ABABACAD", x"AFB1B2B2",
									 -- x"B0B0B0B1", x"B0B1B5BA", x"BAB9BBBF", x"C2C2C2C3", x"C6C5C5C8", x"C9C7C5C6", x"C8C9C8C6", x"C5C6C6C4",
									 -- x"C4C4C4C4", x"C4C2BFBD", x"BAB9B7B4", x"B4B5B3AF", x"AEA9AAA9", x"A4A1A3A3", x"A3A3A3A0", x"9D9C9C9E",
									 -- x"85888B8D", x"8E909395", x"989EA2A3", x"A2A2A2A1", x"A4A4A5A6", x"A7A7A7A6", x"A4A5A6A7", x"A8A7A4A2",
									 -- x"AAA7A7A8", x"A9A7A5A5", x"A5A5A6A5", x"A5A5A7A8", x"A7A8A9A8", x"A8A8A9AB", x"ABACACAB", x"ABACABA9",
									 -- x"ACAAA7A2", x"A1A4A6A6", x"A5A4A3A3", x"A3A3A1A0", x"9E9D9B9A", x"99979391", x"93929190", x"91919090",
									 -- x"908D8B8A", x"87858486", x"87878787", x"86858381", x"85858481", x"8080807E", x"7B787677", x"77777779",
									 -- x"76767678", x"79797775", x"7A797879", x"7977787A", x"7A7C7B7C", x"807F7D7E", x"82848484", x"84878888",
									 -- x"8C8C8D8F", x"8F909397", x"96989C9E", x"A0A2A5A6", x"A7A7A9AC", x"AEAFB1B4", x"B3B5B9BB", x"BCBEC0C1",
									 -- x"C2C3C3C2", x"C1C2C1BF", x"BCBCBCBC", x"BBBAB9B9", x"BBBABABA", x"BABABABA", x"BAB9B9B9", x"BABBBBBB",
									 -- x"BDBDBDBD", x"BBBBBCBE", x"C1C1C0BF", x"BEBFC2C4", x"C5C4C4C6", x"C7C6C7C9", x"CBCDCFD0", x"D1D2D3D4",
									 -- x"D4D5D5D3", x"D2D1CFCD", x"CBCACAC8", x"C6C4C4C3", x"C3C0BFC0", x"C0BDBCBC", x"BBBABBBB", x"BAB7B7BA",
									 -- x"B8B7B6B6", x"B7B8B9B9", x"BDC1C3C7", x"C9C7C8D0", x"CCCDCFD0", x"D2D3D4D4", x"D9D9DADA", x"DAD9D9D8",
									 -- x"D9D9DAD9", x"D9DADBDC", x"DBDBDCDD", x"DEDEDDDD", x"DDDEDFE0", x"E2E2E2E1", x"E2E3E2E0", x"E0E1E2E0",
									 -- x"DFDFDDDD", x"DEE1E0DE", x"DDDDDDDE", x"DFDEDDDC", x"DCD8D6D6", x"D4D0CFD1", x"CCCAC9CA", x"C9C4C0BE",
									 -- x"BAB9B7B7", x"B7B5B1AE", x"ABA8A8A8", x"A19C9A97", x"9695918E", x"8D8C8883", x"87858381", x"7F7D7C7C",
									 -- x"7E7B7775", x"72706D6B", x"6A686563", x"63636261", x"5C605E61", x"5F5A5C59", x"5A575556", x"57565657",
									 -- x"58565557", x"57555456", x"5A5A5957", x"585A5A58", x"54575A5F", x"605B595C", x"61616161", x"62646566",
									 -- x"656A676A", x"6B666A6D", x"6B6E6E6A", x"6A6D6F6E", x"70717174", x"78777880", x"7D7F7D7C", x"7F7F7E81",
									 -- x"868A8A8A", x"8E8F8D8E", x"91919294", x"97989795", x"93969898", x"9BA1A4A2", x"A1A2A3A4", x"A5A7A9AB",
									 -- x"AAAAA9A8", x"A8A9ACAF", x"B1B0AEAE", x"B3B5B0A7", x"A9ABACAA", x"AAACACAB", x"AEAFAFB1", x"B3B5B6B5",
									 -- x"B1B2B3B6", x"B7B7BABE", x"B9BABDC2", x"C5C4C3C2", x"C7C6C7CA", x"CCCAC9CA", x"C8C9C9C7", x"C7C8C7C5",
									 -- x"C8C7C7C7", x"C6C5C3C1", x"BABAB9B6", x"B4B4B2AF", x"AFAAA9A8", x"A3A2A4A5", x"A3A2A1A0", x"9F9D9B99",
									 -- x"7E808487", x"8A8E9396", x"999EA2A2", x"A0A0A2A2", x"A2A3A4A6", x"A7A7A6A5", x"A2A4A5A5", x"A5A4A3A3",
									 -- x"AAA7A5A6", x"A8A7A4A3", x"A7A7A7A6", x"A5A5A6A7", x"A4A7A9A9", x"A7A7A8AA", x"ACABA9A8", x"A9ABAAA8",
									 -- x"A6A7A7A5", x"A4A4A3A1", x"A3A2A2A2", x"A1A1A09F", x"9D9C9B99", x"97959392", x"91908E8E", x"8F8F8F8F",
									 -- x"908E8C8A", x"87858587", x"88888886", x"85848484", x"8383817F", x"7F807F7D", x"7A787777", x"77757575",
									 -- x"75747577", x"79797673", x"77767677", x"77757678", x"797C7C7B", x"7D7D7C80", x"82848584", x"85888989",
									 -- x"8E8E8F90", x"90919498", x"97999C9F", x"A0A2A5A7", x"A7A7A9AC", x"AFB0B1B3", x"B2B5B9BC", x"BDBFC0C2",
									 -- x"BFC0C1C0", x"C0C0C0BE", x"BEBEBEBD", x"BCBBBAB9", x"B9BABABA", x"BABBBBBB", x"BBBAB9B9", x"BABBBCBC",
									 -- x"BDBFBFBE", x"BDBDBEBF", x"C2C2C0BF", x"BFC0C3C4", x"C4C4C5C7", x"C8C7C7C8", x"CBCCCECF", x"D0D0D1D2",
									 -- x"D4D3D3D4", x"D3D0CECE", x"CCCBCAC8", x"C6C5C4C3", x"C2C0C0C0", x"C0BFBDBD", x"BDBCBCBB", x"B9B7B9BD",
									 -- x"BEBEBEBE", x"C0C1C2C2", x"C2C1C2C7", x"CAC5C6CE", x"CBCDCFD1", x"D2D3D5D6", x"D9D9DADB", x"DBDBDAD9",
									 -- x"DCDCDCDB", x"DBDBDBDC", x"DDDCDBDD", x"DFDFDEDC", x"DDDEE0E2", x"E4E5E4E3", x"E1E2E2E0", x"E0E0E0DE",
									 -- x"E1E1DFDE", x"DFE0E0DE", x"DFDEDDDD", x"DEDFDFDF", x"DCDAD7D4", x"D3D3D2D1", x"CECCCBCC", x"CAC6C2C0",
									 -- x"BDBBB9B8", x"B8B5B1AE", x"ABA9ABA8", x"9F9A9B9A", x"97969490", x"8D8C8987", x"88868380", x"7D7C7B7B",
									 -- x"7C797573", x"73726E6A", x"66666563", x"62616060", x"5A5E5D60", x"5F5A5B58", x"5E585353", x"56575655",
									 -- x"56555453", x"52525355", x"59575555", x"585A5956", x"5454595E", x"5B595B5E", x"61616262", x"63636464",
									 -- x"65696568", x"6A66696B", x"666A6C6B", x"6B6E6F6D", x"6F727171", x"75787A7F", x"82827E7D", x"82848386",
									 -- x"8387898D", x"92908E90", x"94949597", x"98989593", x"97999B9A", x"9DA2A4A3", x"A2A3A5A7", x"A8A9AAAB",
									 -- x"AEACA9A8", x"A9ACB0B3", x"B2B3B3B2", x"B1B1B1B1", x"AEAFAEAD", x"ADAFB0AE", x"B1B1B2B4", x"B6B7B7B7",
									 -- x"B4B4B6BA", x"BCBCBDBE", x"BDBEC0C5", x"C7C7C6C6", x"C7C7C8CB", x"CCCBCACA", x"C9CACBCA", x"CAC9C8C6",
									 -- x"C5C4C4C3", x"C3C1C0BE", x"B8B9B8B6", x"B5B4B3B2", x"AFAAA8A8", x"A5A5A6A4", x"A4A2A0A1", x"A29F9A96",
									 -- x"76797D82", x"878C9094", x"959BA1A1", x"9FA0A2A3", x"A2A2A3A5", x"A6A6A4A3", x"A2A3A3A2", x"A1A2A5A8",
									 -- x"A7A6A5A5", x"A6A6A4A3", x"AAA9A9A7", x"A6A6A6A6", x"A4A6A8A9", x"A8A7A7A7", x"A9A9A7A6", x"A7A9A9A7",
									 -- x"A3A5A6A5", x"A5A4A3A0", x"A2A1A0A0", x"A09F9E9D", x"9B9B9A97", x"95939394", x"908F8E8E", x"8E8F8F8F",
									 -- x"8E8E8C8A", x"87858585", x"88888786", x"83838486", x"7F807F7F", x"80817D79", x"7C7A7877", x"76757473",
									 -- x"75757577", x"78787675", x"73737476", x"76757678", x"797C7B7A", x"7D7E7E81", x"82848585", x"86898B8B",
									 -- x"8E8F9090", x"91929497", x"989A9C9E", x"9FA0A2A4", x"A8A7A9AD", x"AFAFB0B1", x"B3B6BABD", x"BEBFC0C1",
									 -- x"BEBFC0BF", x"BFC0BFBD", x"BEBEBEBE", x"BDBDBCBC", x"BBBBBBBB", x"BBBBBBBB", x"B9B9B8B9", x"BABCBEBF",
									 -- x"BEC0C2C1", x"BFC0C0C0", x"C0C0C1C2", x"C2C3C4C4", x"C4C4C5C6", x"C7C7C7C8", x"C9CACCCD", x"CFD0D2D3",
									 -- x"D4D1D1D4", x"D3CFCED0", x"CDCCCAC8", x"C6C5C4C3", x"C2C1C1C1", x"C1C0BFBE", x"BFBFBFBD", x"BBBABDC0",
									 -- x"BDBEBFC0", x"C2C2C2C1", x"C2C3C4C7", x"CAC7C6CB", x"CACDD1D3", x"D3D4D7D9", x"D8D9D9DA", x"DBDCDDDD",
									 -- x"DEDEDEDD", x"DCDCDCDC", x"DEDEDDDE", x"E0E1E0E0", x"E1E1E2E4", x"E5E5E4E3", x"E2E2E3E2", x"E1E1E0DE",
									 -- x"E2E2E1DF", x"DFE0DEDC", x"DFDEDDDD", x"DEDFE0E0", x"DCDBD7D3", x"D3D5D4D0", x"D2CFCCC9", x"C8C6C4C3",
									 -- x"BFBDBAB8", x"B7B5B2B0", x"ABA9A9A7", x"A09B9D9D", x"99979591", x"8E8D8C8C", x"8987837F", x"7D7B7B7B",
									 -- x"78757271", x"71706C69", x"64646362", x"61616161", x"5C5E5A5C", x"5B585C5A", x"5D595656", x"58585553",
									 -- x"55565653", x"51525353", x"55545253", x"56585654", x"5754595D", x"59595D5C", x"60616161", x"62626364",
									 -- x"64676266", x"6966686A", x"62676B6E", x"7072716F", x"6E747472", x"757B7F84", x"84858180", x"84868587",
									 -- x"8385888D", x"928F8D92", x"95969798", x"99999795", x"9B9D9E9D", x"9EA1A2A1", x"A3A5A7A9", x"AAACADAE",
									 -- x"B2B0AEAD", x"AEB1B3B5", x"B5B6B6B5", x"B1B0B5BB", x"B4B3B1AF", x"B0B2B3B2", x"B5B4B4B6", x"B8B9BABB",
									 -- x"BBBABBBE", x"BFBFBEBF", x"C5C4C4C6", x"C8C8C9CB", x"C9C9CACB", x"CCCBCAC9", x"CACBCCCC", x"CBCAC8C6",
									 -- x"C6C5C5C5", x"C4C3C0BF", x"BAB8B6B5", x"B5B5B3B1", x"AEA9A8A9", x"A8A7A6A1", x"A5A3A2A2", x"A2A09B97",
									 -- x"777A7E82", x"868A8D8F", x"93999FA1", x"A0A1A2A3", x"A3A3A4A5", x"A5A5A4A2", x"A0A1A2A1", x"9FA0A4A7",
									 -- x"A3A5A6A5", x"A4A4A5A6", x"A7A7A6A5", x"A5A5A4A4", x"A6A5A6A7", x"A8A7A5A4", x"A5A7A8A6", x"A5A6A6A6",
									 -- x"A5A4A29E", x"9EA1A3A4", x"A1A09F9F", x"9F9E9D9C", x"97979593", x"91909192", x"8F8E8D8D", x"8E8E8E8E",
									 -- x"8B8C8B89", x"87858483", x"87878583", x"81808183", x"8181807F", x"7F7E7A76", x"7B797776", x"76767676",
									 -- x"74767676", x"75747576", x"74747577", x"77767779", x"797B797A", x"7F808082", x"82848686", x"888B8C8C",
									 -- x"8E909191", x"92949799", x"989A9C9D", x"9E9FA1A3", x"A7A7A9AC", x"AEAEAFB1", x"B5B8BBBE", x"BEBFBFC0",
									 -- x"C0C2C2C1", x"C1C1C1BF", x"BEBEBEBE", x"BEBEBDBD", x"BDBDBEBE", x"BEBDBDBD", x"B9B9B9B9", x"BABCBEBF",
									 -- x"BEC1C2C1", x"C0C1C2C1", x"BFBFC0C1", x"C2C3C3C3", x"C4C5C5C5", x"C6C7C8C8", x"C8CACBCD", x"CED0D2D3",
									 -- x"D3D1D1D3", x"D2CFCED0", x"CDCCC9C7", x"C6C6C4C4", x"C4C3C3C2", x"C2C2C0BF", x"C0C1C2C0", x"BEBEBFC1",
									 -- x"BDBDBFC1", x"C2C2C1BF", x"C0C7C8C6", x"C9CBC9C9", x"CBCED2D3", x"D4D5D8DA", x"DBDADADA", x"DBDDDEE0",
									 -- x"E0E0E0DF", x"DEDDDDDD", x"DEDFE0E0", x"E0E1E2E3", x"E4E4E3E4", x"E5E5E4E4", x"E4E4E4E5", x"E4E2E1E0",
									 -- x"E0E2E2E1", x"E0E1DFDC", x"DEDDDDDE", x"DFE0E0E0", x"DDDCD9D4", x"D4D6D5D0", x"D0CECBC9", x"C8C7C5C3",
									 -- x"C0BEBAB8", x"B6B5B3B2", x"ADA8A7A6", x"A19E9E9D", x"9996938F", x"8B898B8C", x"8C898580", x"7C7A7878",
									 -- x"78757370", x"6E6B6866", x"65625F5E", x"5F5F605F", x"5C5D5859", x"59575B5A", x"59585756", x"56555351",
									 -- x"54565553", x"52525251", x"52525354", x"55555555", x"55525960", x"5E5E5E58", x"60606161", x"61626465",
									 -- x"64676266", x"69676A6C", x"66696D70", x"72747473", x"70787975", x"777D848A", x"84868482", x"84848385",
									 -- x"8A8B8B8E", x"918E8E94", x"94949698", x"9A9C9D9D", x"9A9D9FA0", x"A2A4A4A4", x"A6A7A9AB", x"ADAEB0B1",
									 -- x"B3B2B2B3", x"B4B5B5B5", x"BCB8B6B8", x"BBBBBBBB", x"B8B6B3B0", x"B2B6B8B8", x"BCB9B8BA", x"BBBCBDC0",
									 -- x"C2C0BFC1", x"C3C2C3C4", x"C9C7C7C8", x"C9C9CACC", x"CBCBCCCC", x"CDCECDCC", x"CBCBCCCC", x"CBC8C6C5",
									 -- x"C5C5C5C5", x"C4C2BFBC", x"BFBAB5B3", x"B4B3AFAC", x"AEA8A7A7", x"A6A7A6A1", x"A2A2A2A1", x"A09D9B99",
									 -- x"77797C81", x"85898C8D", x"94999EA0", x"A0A1A1A0", x"A0A0A0A0", x"A1A1A09F", x"9D9FA1A0", x"9F9FA0A1",
									 -- x"A0A3A5A4", x"A2A4A6A8", x"A4A4A4A4", x"A5A5A5A4", x"A6A4A3A4", x"A6A6A4A1", x"A2A6A7A6", x"A4A3A3A3",
									 -- x"A1A19F9D", x"9D9FA0A0", x"A09F9E9E", x"9D9C9B9A", x"95949290", x"8F8F8F8F", x"8D8C8C8C", x"8C8C8C8B",
									 -- x"8C8D8D8B", x"88888785", x"88878683", x"81808080", x"81817F7D", x"7D7E7D7B", x"7C7B7976", x"75767675",
									 -- x"74767775", x"72727476", x"75757577", x"76757678", x"787A7879", x"7F818183", x"81848787", x"898C8E8E",
									 -- x"8E909293", x"94979A9C", x"999A9C9E", x"9FA0A3A5", x"A5A6A9AC", x"AEAEB1B4", x"B7BABCBE", x"BEBEBFC0",
									 -- x"C1C2C3C2", x"C2C2C2C0", x"C0C0C0BF", x"BFBEBDBD", x"BCBDBDBE", x"BEBEBDBD", x"BBBBBBBB", x"BABBBCBE",
									 -- x"BDC1C2BF", x"BFC1C2C1", x"C3C1BFBE", x"BFC1C2C3", x"C5C6C6C5", x"C6C7C8C8", x"CACBCCCD", x"CECFD1D2",
									 -- x"D2D1D1D2", x"D1CFCECF", x"CECBC9C7", x"C7C7C5C4", x"C5C5C4C3", x"C3C4C2C0", x"C1C2C2C1", x"C0C1C1C1",
									 -- x"C2C3C4C5", x"C6C6C5C4", x"C1CBCCC8", x"CBCECDCC", x"CED0D2D3", x"D4D5D8DA", x"DEDEDDDC", x"DCDEDFE0",
									 -- x"E1E2E2E1", x"E0DFDFDF", x"DDDFE1E2", x"E1E0E2E3", x"E4E3E3E3", x"E4E5E5E4", x"E2E2E2E3", x"E3E1E0E0",
									 -- x"DFE1E2E2", x"E2E2E1DF", x"DEDEDFE0", x"E1E1E0DF", x"DEDDDBD7", x"D6D6D4D1", x"CCCCCCCB", x"CAC9C6C2",
									 -- x"C1BEBBB8", x"B5B4B2B1", x"AFA8A5A5", x"A19F9F9C", x"9B97938F", x"8B88888A", x"89878480", x"7D7A7978",
									 -- x"7574716F", x"6D6B6867", x"6764605E", x"5E5E5E5D", x"5A5B5759", x"59575A57", x"58595854", x"52525353",
									 -- x"52515152", x"5251504F", x"50525456", x"55535456", x"5653555A", x"5C5F5F5C", x"5F606161", x"60626467",
									 -- x"62666265", x"6865696C", x"6D6D6D6D", x"6F727373", x"737A7B77", x"797D838A", x"87898886", x"88868487",
									 -- x"8C8E8E8E", x"91929399", x"9797999A", x"9C9D9E9F", x"9E9FA1A3", x"A5A6A6A6", x"A8A9ACAD", x"AFB0B2B3",
									 -- x"B1B2B4B6", x"B8B8B8B8", x"B9BABBBD", x"BFBEBDBB", x"B8B8B6B4", x"B6BABDBE", x"BEBBB9BC", x"BDBDBEC1",
									 -- x"C3C1C1C2", x"C3C4C6C8", x"C8C7C8CB", x"CCCBC9C9", x"CACBCBCB", x"CCCECFCE", x"CDCCCBCB", x"C9C7C5C6",
									 -- x"C4C4C4C3", x"C2BFBCB9", x"BBB6B2B3", x"B4B2AEAB", x"AEA8A5A2", x"A1A4A6A2", x"9FA0A1A0", x"9C999899",
									 -- x"77787A7E", x"83878B8C", x"93979A9B", x"9D9F9F9D", x"9B9B9A9A", x"9B9B9B9B", x"999A9C9D", x"9C9C9C9D",
									 -- x"9FA2A3A2", x"A1A4A6A6", x"A5A5A4A5", x"A6A6A5A4", x"A3A2A0A1", x"A2A2A2A1", x"A2A4A4A3", x"A3A3A3A1",
									 -- x"9C9FA0A0", x"9F9F9C9A", x"9E9D9C9C", x"9C9B9998", x"97949290", x"8F8F8E8D", x"8C8B8C8C", x"8C8B8A89",
									 -- x"8C8D8C89", x"88888988", x"87868584", x"83828180", x"7E7F7F7D", x"7E80807F", x"7D7D7A77", x"75767472",
									 -- x"77777876", x"74737475", x"75747575", x"75747578", x"7679797A", x"7E7F8084", x"81848788", x"8A8D8F8F",
									 -- x"8E919393", x"94989B9B", x"9A9B9D9E", x"9FA1A3A6", x"A5A7ABAD", x"ADAEB2B7", x"B9BBBDBE", x"BEBEBFC0",
									 -- x"C0C2C3C2", x"C2C3C3C2", x"C2C2C1C1", x"C0BFBEBD", x"BDBDBEBE", x"BDBCBBBB", x"BDBDBDBD", x"BCBCBDBE",
									 -- x"BEC2C2BF", x"BFC2C3C2", x"C4C2C0C0", x"C1C3C4C4", x"C5C7C8C7", x"C7C9C9C8", x"CACBCCCC", x"CDCECFD1",
									 -- x"D1D2D2D0", x"CFD0CFCE", x"CECBC8C7", x"C7C7C6C5", x"C5C6C6C4", x"C5C6C5C3", x"C4C4C3C1", x"C2C4C4C2",
									 -- x"C4C4C4C4", x"C5C6C6C6", x"C7CECFCC", x"CED0D1D3", x"D3D3D3D4", x"D6D8D9DB", x"E0E0E0E0", x"E0E0E1E1",
									 -- x"E3E3E4E4", x"E3E2E1E1", x"E0E1E2E3", x"E3E2E2E2", x"E3E2E3E3", x"E4E4E3E3", x"E2E0E1E2", x"E2E0DFE0",
									 -- x"E2E3E3E2", x"E2E3E3E2", x"DFDFE0E2", x"E3E2E1E0", x"DFDFDDDB", x"D8D6D4D3", x"CDCECECC", x"CCCAC6C1",
									 -- x"C0BEBCB9", x"B5B3B0AF", x"ADA7A5A5", x"A1A09F9C", x"9D999592", x"8F8A8889", x"84838280", x"7E7B7978",
									 -- x"74716D6C", x"6C6B6866", x"6564615F", x"5D5C5C5C", x"585A5659", x"59575955", x"595A5854", x"52525454",
									 -- x"504C4B4F", x"52504F4F", x"4F505355", x"54515154", x"57565251", x"565B5D60", x"5C5E6060", x"60606264",
									 -- x"61666265", x"6764696D", x"716F6E6E", x"6F717272", x"787B7A79", x"7C7F8389", x"8B8C8A89", x"8C8C8A8B",
									 -- x"8A8F9090", x"9496989C", x"9B9C9D9E", x"9D9D9D9D", x"A2A2A3A4", x"A5A6A6A7", x"AAACAEB0", x"B1B2B2B3",
									 -- x"B1B4B6B8", x"B9BABBBC", x"B6BCC0BF", x"BDBDBDBB", x"BABBBBB9", x"BABDBFC0", x"BEBBBBBE", x"BFBEBEC0",
									 -- x"C3C2C2C2", x"C3C4C7CB", x"C9C8CACD", x"CECDCBCB", x"CACBCAC9", x"CBCECFCE", x"CECCCACA", x"C8C6C6C7",
									 -- x"C9C8C6C4", x"C3C0BEBC", x"B5B3B3B5", x"B4B0ACAB", x"ABA7A4A1", x"9FA2A49F", x"9E9FA09F", x"9B979696",
									 -- x"7C7C7C7E", x"81858889", x"92949597", x"9A9D9D9C", x"9A999898", x"999A9B9A", x"97979797", x"98999B9D",
									 -- x"9FA1A1A0", x"A1A4A6A4", x"A6A5A5A5", x"A5A5A3A2", x"A0A09F9F", x"9F9FA1A2", x"A1A1A1A1", x"A3A5A4A2",
									 -- x"A1A1A09D", x"9C9D9D9C", x"9D9C9B9B", x"9A999897", x"9794918F", x"8F8E8D8B", x"8C8C8C8D", x"8D8C8A88",
									 -- x"8A8A8985", x"83858786", x"83828182", x"83838280", x"7D808281", x"80807E7D", x"78797977", x"77787674",
									 -- x"79797979", x"78777574", x"76757577", x"7777797B", x"74797B7B", x"7D7D7E84", x"81858789", x"8B8E8F8F",
									 -- x"8F929493", x"93969898", x"9B9C9D9E", x"9E9FA2A4", x"A7AAADAF", x"ADADB1B7", x"B9BBBDBE", x"BEBEBFC1",
									 -- x"C2C4C5C4", x"C5C6C6C5", x"C3C2C2C2", x"C1C0BFBF", x"C0C0C0C0", x"BEBDBBBA", x"BCBDBEBE", x"BEBDBEC0",
									 -- x"C0C4C4C0", x"C0C3C5C4", x"C3C3C3C4", x"C6C7C7C6", x"C5C8C9C9", x"C9CBCAC7", x"C9CACBCB", x"CCCDCFD1",
									 -- x"D1D3D2CF", x"CED0CFCD", x"CECBC8C7", x"C7C8C7C6", x"C5C6C6C5", x"C5C7C7C4", x"C8C7C4C2", x"C4C7C6C4",
									 -- x"C9C8C6C6", x"C7C9CBCC", x"CCD0D0D0", x"D0CFD2D9", x"D7D6D5D6", x"D8DADCDC", x"E0E0E1E2", x"E3E3E3E3",
									 -- x"E4E4E5E5", x"E5E4E3E4", x"E4E4E3E5", x"E6E5E3E1", x"E2E2E3E4", x"E4E3E1E0", x"E4E2E3E4", x"E4E2E2E3",
									 -- x"E6E7E5E2", x"E1E2E3E3", x"E1E1E2E3", x"E3E3E2E1", x"E1E0DFDD", x"DAD6D4D4", x"D3D3D0CC", x"CAC9C6C2",
									 -- x"BFBFBDBA", x"B6B2AEAC", x"AAA5A4A5", x"A1A0A19F", x"9B989594", x"918C8988", x"85848380", x"7D797673",
									 -- x"77726B69", x"6A69645F", x"5F60605E", x"5A59595B", x"595A5557", x"57565956", x"56585754", x"53535251",
									 -- x"4F49484E", x"52504F51", x"4D4E5053", x"524F4F51", x"52575452", x"5758585C", x"595B5E5F", x"5E5E5F61",
									 -- x"62686567", x"69666B70", x"72727274", x"75757473", x"7E7E7B7C", x"8285878C", x"8D8C8888", x"8E8F8D8D",
									 -- x"8D959694", x"9699999A", x"9A9C9E9F", x"9F9F9E9D", x"A1A0A0A2", x"A3A5A8AA", x"ABADB1B3", x"B3B3B2B1",
									 -- x"B5B7B9BA", x"B9BBBDC0", x"C0C0BDBB", x"BFC4C1B9", x"BCBEBFBE", x"BDBEBFBF", x"C0BDBEC2", x"C3C0BFC2",
									 -- x"C5C5C5C5", x"C5C5C9CE", x"CCCACACD", x"CECECFD0", x"CECECDCB", x"CCCFD1CF", x"CFCBC9C9", x"C8C6C7C9",
									 -- x"C8C5C2BF", x"BDBCBAB9", x"B5B6B8B8", x"B3ABA6A5", x"A7A5A5A4", x"A0A2A19B", x"9FA0A19F", x"9C989594",
									 -- x"7B7B797C", x"8284858A", x"91929393", x"93939596", x"98969494", x"95969695", x"96979694", x"95999B9B",
									 -- x"9C9D9FA0", x"A1A2A4A5", x"A5A5A4A3", x"A5A6A4A0", x"A2A2A09F", x"9E9F9FA0", x"A2A3A19E", x"9EA0A09F",
									 -- x"A09F9F9F", x"9E9D9A97", x"9C9D9D9B", x"9A9A9996", x"9895908C", x"8E918F8B", x"8B8A8A8A", x"8B8A8988",
									 -- x"85868583", x"83858583", x"82838484", x"84858583", x"827F7F81", x"817D7A7B", x"77787876", x"77797977",
									 -- x"7778797A", x"79767472", x"77767574", x"76797A78", x"767B7A78", x"7B7D7D7F", x"84818389", x"8C8D8D90",
									 -- x"8F909292", x"9192979C", x"9C9D9E9E", x"9E9FA2A4", x"A8ABAFB1", x"AFAEB2B7", x"BABCBEBF", x"BFBFC1C2",
									 -- x"C5C5C4C4", x"C4C4C4C4", x"C3C3C4C3", x"C2C2C3C3", x"C2C3C2C1", x"BFBFC0C2", x"C0BFBEBE", x"BEBEBCBA",
									 -- x"BFC0C0BF", x"BFC2C4C5", x"C5C6C5C5", x"C5C5C6C7", x"C7C8C9C9", x"C8C8C9CA", x"CCCCCCCC", x"CDCED1D3",
									 -- x"D3D3D3D2", x"D1D0D0D0", x"CDCBC8C7", x"C8C8C8C8", x"C4C5C7C9", x"CAC9C8C6", x"C8C8C8C7", x"C6C7C9CA",
									 -- x"CACAC9CA", x"CACBCCCD", x"D1D2D3D4", x"D4D4D5D5", x"D5D7DADB", x"DADBDEE1", x"E4E3E3E5", x"E6E5E5E8",
									 -- x"E7E7E8E8", x"E8E8E7E7", x"E8E8E7E6", x"E6E5E4E4", x"E4E4E3E3", x"E4E4E3E2", x"E1E2E3E4", x"E5E5E5E4",
									 -- x"E6E6E6E5", x"E5E5E5E5", x"E5E4E3E2", x"E1E2E3E3", x"E3E0DFDE", x"DAD8D7D3", x"D4D4D2CD", x"CAC9C7C4",
									 -- x"C2BFBCB9", x"B5B1AFB0", x"ACAAA7A5", x"A4A29F9C", x"9B959294", x"928D8989", x"8B838082", x"7D787674",
									 -- x"6F6D6A68", x"67666360", x"6060605E", x"5B59595B", x"58565252", x"53555555", x"56565553", x"54555450",
									 -- x"4F49474A", x"4C4B4A4D", x"48494C4F", x"4E4B4F55", x"54565452", x"5253555B", x"5A5E5E5D", x"5E5D5C5D",
									 -- x"64666867", x"64656A6F", x"736F6F73", x"7372767D", x"807C7E83", x"8382878F", x"8E8B8A8E", x"918F8C8B",
									 -- x"90949695", x"94989A9A", x"9A9DA1A3", x"A3A2A2A2", x"A3A2A2A5", x"A9ABACAB", x"A8B0B2AF", x"B2B4B4B5",
									 -- x"B4B8BBBC", x"BEC1C1C1", x"BEBFC2C5", x"C6C3C3C4", x"C5C0BCBC", x"BDBEC1C4", x"C0C1C3C4", x"C2BFBFC2",
									 -- x"C9C6C5C6", x"C7C8C9CC", x"CBCDD0D1", x"D1D0CFCE", x"D2CECDD0", x"D0CECED1", x"CECDCCCC", x"CECDCAC7",
									 -- x"C4C4C1BB", x"BABCBCB9", x"B9B5B2B0", x"ADAAABAE", x"A8A8A6A3", x"A2A2A09E", x"A2A29E9B", x"9B979191",
									 -- x"7B7B7A7C", x"8283858A", x"8E8F9191", x"91929394", x"93949596", x"9694918E", x"93959594", x"95979897",
									 -- x"999B9C9E", x"9E9FA0A1", x"A2A3A3A3", x"A4A5A3A0", x"A1A0A0A0", x"A1A1A2A2", x"A1A2A19F", x"9EA0A0A0",
									 -- x"9F9E9D9C", x"9C9C9B99", x"9B9A9896", x"96979592", x"9193928E", x"8C8C8C8B", x"8C8B8B8A", x"89888787",
									 -- x"83848382", x"82838381", x"81828281", x"83858482", x"807F7F81", x"817E7C7B", x"7B7B7A77", x"78797977",
									 -- x"78797A7A", x"7A787574", x"76767574", x"75787775", x"777B7B79", x"7C7E7E80", x"82828387", x"8B8D8F90",
									 -- x"8F929595", x"9494979B", x"9C9D9E9F", x"A0A1A3A5", x"A6A8ACAF", x"AFAFB2B7", x"BABDC1C3", x"C3C2C2C3",
									 -- x"C9C9C8C7", x"C6C5C4C4", x"C4C5C5C5", x"C4C2C2C2", x"C2C3C3C3", x"C1C1C1C1", x"C0C0C0C0", x"C0C0BFBE",
									 -- x"C0C1C2C1", x"C1C4C5C6", x"C7C7C7C7", x"C7C7C8C9", x"C9CACBCA", x"C9C8C9CA", x"CBCCCCCD", x"CECFD2D4",
									 -- x"D3D4D4D3", x"D2D1D0CF", x"CCCBC9C8", x"C8C8C7C7", x"C5C6C7C9", x"CACAC9C9", x"C9C9C9C8", x"C8C8C9CA",
									 -- x"CBCBCCCD", x"CECFD0D1", x"D3D4D5D6", x"D6D6D7D8", x"D8DADCDD", x"DCDEE1E5", x"E4E3E5E8", x"E8E7E7E9",
									 -- x"E9EAEAEA", x"EAEAEAEA", x"EAEAE9E8", x"E7E7E6E6", x"E6E5E4E4", x"E5E5E4E3", x"E2E3E3E3", x"E4E5E5E6",
									 -- x"E4E5E6E7", x"E7E6E4E3", x"E6E5E4E3", x"E3E3E3E4", x"E2DFDFDF", x"DBDAD9D5", x"D2D2D1CE", x"CCCCCAC8",
									 -- x"C3C0BDBB", x"B8B3B1B1", x"ABACACA8", x"A29E9C9D", x"9E989494", x"938E8B8B", x"867F7E80", x"7C797876",
									 -- x"6E6B6867", x"66656260", x"5C5D5C5A", x"57555657", x"55545353", x"55555453", x"53545452", x"5253514F",
									 -- x"4E4C4D4E", x"4B47494E", x"49494B4C", x"4C4C4D50", x"4E525251", x"5253555B", x"5A5D5C5B", x"5D5C5B5D",
									 -- x"60646767", x"66686C71", x"73717276", x"77777B80", x"80808182", x"83858A8F", x"8D8D8F94", x"96959392",
									 -- x"90959796", x"979A9C9B", x"9B9DA0A0", x"9FA0A4A8", x"A6A5A5A7", x"AAADAEAF", x"AEB4B4B2", x"B5B8B7B6",
									 -- x"B8BCBEBE", x"BEC0C1C2", x"C4C2C3C4", x"C5C4C5C7", x"C4C0BEC0", x"C1C1C2C4", x"C3C3C4C5", x"C4C2C4C7",
									 -- x"C7C5C6C8", x"CACACCCD", x"CFD0D1D1", x"D1D0CFCE", x"CED1D0CC", x"CDD1D0CC", x"CCCCCDCD", x"CCCAC7C6",
									 -- x"C2C2C0BD", x"BCBDBCBA", x"B9B5B0AD", x"ABAAACAF", x"A8A8A6A4", x"A2A2A09E", x"9C9C9895", x"97959192",
									 -- x"7A7C7B7D", x"81828489", x"8A8C8E90", x"90909192", x"95949292", x"91919090", x"91939494", x"95969694",
									 -- x"999A9C9D", x"9E9E9F9F", x"9FA1A3A3", x"A3A3A19E", x"A0A0A0A1", x"A1A2A2A3", x"9EA0A09F", x"9D9E9F9F",
									 -- x"9E9C9B9A", x"9A9B9B9B", x"9B999594", x"95979591", x"8F908F8C", x"8A898989", x"8B8B8B8A", x"87868686",
									 -- x"83848483", x"83838280", x"81817F7E", x"81838381", x"80818181", x"80807D7A", x"7C7C7A78", x"78797877",
									 -- x"7778797A", x"79787674", x"74757474", x"76787775", x"787C7C7B", x"7E7F7F81", x"82838486", x"8A8E9090",
									 -- x"92949796", x"9596999B", x"9E9E9FA0", x"A1A2A3A5", x"A5A7AAAE", x"B0B2B5B9", x"BDBFC3C5", x"C5C5C5C6",
									 -- x"CCCCCBCA", x"C8C7C5C5", x"C5C6C7C6", x"C5C4C3C3", x"C3C4C5C5", x"C4C3C2C1", x"C1C1C2C2", x"C1C0C0C0",
									 -- x"C0C2C3C2", x"C3C5C6C6", x"C7C8C8C8", x"C8C9CACB", x"CBCBCCCB", x"CBCBCBCC", x"CDCDCECE", x"CED0D1D3",
									 -- x"D3D3D4D5", x"D4D2D0CF", x"CCCBC9C8", x"C8C8C6C5", x"C6C6C7C9", x"CACBCCCC", x"CDCDCDCD", x"CDCDCDCE",
									 -- x"CDCED0D1", x"D2D3D4D5", x"D7D8D9DA", x"DADBDBDC", x"DCDEDFDF", x"DEE0E3E6", x"E5E5E8EB", x"ECEBEAEA",
									 -- x"ECECECED", x"EDEDEDEC", x"EDECECEB", x"EAE9E9E8", x"E7E7E6E6", x"E6E6E5E5", x"E5E4E4E3", x"E4E5E6E7",
									 -- x"E5E6E7E7", x"E7E6E5E4", x"E6E6E5E4", x"E4E4E4E4", x"E3E0E0E0", x"DCDBDAD6", x"D7D6D3D0", x"CDCCC9C6",
									 -- x"C4C1BFBE", x"BBB7B3B2", x"ADAEAEAA", x"A49F9C9C", x"A09B9696", x"94908C8C", x"86807F7F", x"79757472",
									 -- x"6D6B6866", x"6564605E", x"5C5C5B58", x"56545556", x"55545353", x"54555453", x"51535351", x"5050504F",
									 -- x"4B4B4B4C", x"4945474B", x"4A4B4B4B", x"4D4F4F4E", x"4C515151", x"5455565B", x"5B5E5D5C", x"5E5D5C5F",
									 -- x"62666969", x"67686B6F", x"71737577", x"797B7D7F", x"81858583", x"84898D8E", x"8C8D9296", x"97969595",
									 -- x"92979998", x"999C9E9D", x"9B9EA09F", x"9EA0A5AA", x"ACABABAB", x"ABABACAD", x"AFB2B1B1", x"B6B9B7B6",
									 -- x"B7BBBFC0", x"C1C3C4C5", x"C5C3C2C3", x"C4C4C4C5", x"C5C3C3C4", x"C5C4C3C3", x"C4C4C4C4", x"C3C3C6CA",
									 -- x"C5C5C6C9", x"CBCBCBCD", x"D1D0D0D1", x"D2D2D0CF", x"CED1D1CE", x"CED1CFCB", x"CECFCFCE", x"CCCAC8C7",
									 -- x"C1BEBCBC", x"BCBBBBBB", x"B8B3AEAC", x"ABABACAE", x"A8A8A6A4", x"A2A2A09D", x"9C9B9693", x"94939193",
									 -- x"797D7D7E", x"81828388", x"86898C8E", x"8E8F8F90", x"9593918F", x"8F909293", x"91929394", x"95959595",
									 -- x"999A9C9D", x"9D9D9D9E", x"9EA0A2A1", x"A0A09F9E", x"A0A0A09F", x"9FA0A0A0", x"9D9E9F9E", x"9C9B9C9D",
									 -- x"9C9B9999", x"98999A9A", x"98979594", x"95969593", x"938F8A89", x"8B8C8A88", x"898A8B89", x"87858688",
									 -- x"85848483", x"8383817E", x"82817E7D", x"7F828280", x"83848380", x"7E7F7D79", x"7A797876", x"76777777",
									 -- x"76777878", x"78767574", x"74747474", x"77797978", x"797C7C7B", x"7E7F7F82", x"83868786", x"898F9291",
									 -- x"96989795", x"95989C9F", x"A1A1A2A2", x"A2A2A3A3", x"A7A7AAAF", x"B3B6B9BD", x"C1C2C3C4", x"C4C6C9CA",
									 -- x"CCCBCBCA", x"C9C7C6C6", x"C6C6C7C7", x"C6C5C5C5", x"C4C5C5C5", x"C5C4C3C2", x"C2C3C3C2", x"C0BFBFBF",
									 -- x"C0C2C3C3", x"C4C5C6C5", x"C7C7C8C9", x"C9C9CACB", x"CBCBCCCD", x"CDCECECF", x"CFCFD0CF", x"CFCFCFD0",
									 -- x"D1D2D4D5", x"D5D3D1CF", x"CDCBC8C7", x"C7C6C5C4", x"C6C7C8CA", x"CBCCCECE", x"D0D1D2D2", x"D1D1D1D1",
									 -- x"D0D1D3D3", x"D4D5D7D8", x"DADCDDDE", x"DEDFE0E0", x"E1E2E3E3", x"E2E3E5E6", x"E7E8EAEC", x"EDEDECEC",
									 -- x"EDEDEEEE", x"EFEFEFEF", x"EFEFEEED", x"EDECEBEB", x"E9E8E8E7", x"E7E7E7E7", x"E7E7E6E6", x"E6E7E8E9",
									 -- x"EAE9E7E6", x"E6E7E8E8", x"E7E7E6E6", x"E5E4E4E3", x"E5E2E2E1", x"DDDCDAD6", x"DBD9D6D2", x"CFCCC9C6",
									 -- x"C6C3C0BF", x"BEBAB6B4", x"B2AFABAA", x"A9A6A19C", x"A19C9898", x"96918D8C", x"8883817F", x"7772706F",
									 -- x"6D6B6765", x"64625E5C", x"5C5C5A58", x"55545555", x"5452504F", x"50515354", x"4F50514F", x"4D4C4C4D",
									 -- x"4A484647", x"49494746", x"474B4B4A", x"4C50514E", x"4D515151", x"53545559", x"5A5C5B5C", x"5E5C5B5F",
									 -- x"65686B6A", x"68686C6F", x"72757776", x"797D7F7E", x"85878887", x"888B8D8D", x"8F8F9193", x"94949494",
									 -- x"96999A98", x"999D9F9E", x"9B9DA0A0", x"A0A2A5A8", x"ACADADAD", x"ABABAAAB", x"ABAFAEAF", x"B5B9B8B9",
									 -- x"B7BBC0C3", x"C5C6C5C3", x"C4C4C4C6", x"C6C5C4C2", x"C8C7C8C8", x"C7C5C3C3", x"C5C5C5C4", x"C3C4C7CB",
									 -- x"C7C7C8CB", x"CCCBCCCE", x"D0CFCED0", x"D3D4D3D2", x"D2CECED3", x"D4CFCDD0", x"D0CFCECC", x"CBCAC8C7",
									 -- x"C2BDB9B9", x"B9B7B8BB", x"B5B2AFAE", x"AFAEACAA", x"A9A8A5A2", x"A0A09F9D", x"9E9D9792", x"93918F90",
									 -- x"7A7E7E7D", x"80818286", x"85878B8D", x"8E8E8E8F", x"8F909192", x"92908F8E", x"90909192", x"94949596",
									 -- x"98999A9A", x"9A9A9A9A", x"9C9E9F9E", x"9D9FA09F", x"A1A09F9E", x"9E9E9FA0", x"9E9E9F9E", x"9C9A9A9B",
									 -- x"9A9A9999", x"98979797", x"95959595", x"94929192", x"938F8B8B", x"8E8E8B88", x"898A8B89", x"87868789",
									 -- x"85838282", x"82807D7B", x"83827F7E", x"7F828280", x"8485837E", x"7D7F7E7A", x"7B797776", x"76767777",
									 -- x"77777777", x"77767575", x"75757373", x"75797978", x"797B7B7B", x"7E7E7E82", x"83868888", x"8B919494",
									 -- x"999B9B99", x"989CA1A3", x"A5A5A5A5", x"A5A6A6A5", x"A8A8ABB0", x"B5B9BCBF", x"C3C4C5C6", x"C7C9CCCD",
									 -- x"CDCDCCCB", x"CAC8C7C7", x"C8C8C8C7", x"C7C6C7C7", x"C6C5C5C4", x"C4C4C4C4", x"C2C3C4C3", x"C1BFBFC0",
									 -- x"C0C3C5C5", x"C5C7C7C6", x"C7C8C9C9", x"C9CACBCB", x"CDCDCDCE", x"CFCFD0D0", x"D0D0D1D0", x"CFCFCFCF",
									 -- x"D0D1D2D4", x"D5D4D1CF", x"CDCAC7C5", x"C5C5C5C4", x"C5C7CACC", x"CDCECFD0", x"D0D2D3D3", x"D3D3D3D3",
									 -- x"D4D5D6D5", x"D5D6D8DA", x"DCDDDEE0", x"E0E1E2E3", x"E3E5E7E8", x"E8E8E8E9", x"EBECECEC", x"EDEEEEED",
									 -- x"F0F0F1F1", x"F2F2F2F2", x"F2F1F0F0", x"EEEEEDEC", x"EAEAEAE9", x"E8E8E8E8", x"E9E9E9E9", x"E9EAEAEA",
									 -- x"ECEBEAE9", x"E9E9EAEB", x"E9E9E8E7", x"E6E5E5E4", x"E5E2E3E3", x"DFDDDCD7", x"D9D6D4D3", x"D2D0CECC",
									 -- x"C9C5C1C0", x"BFBBB8B6", x"B5B1ADAC", x"ABA9A49F", x"9F9C9999", x"97928D8A", x"837F7F7D", x"76737270",
									 -- x"6C696664", x"63615E5B", x"5B5B5957", x"55535353", x"504F4D4C", x"4C4D4F4F", x"4C4D4E4D", x"4B49494A",
									 -- x"4A494747", x"494A4846", x"44484A48", x"494C4E4D", x"4C4F4E4E", x"50515256", x"5557585A", x"5C5A585D",
									 -- x"65686B6A", x"696B7075", x"76797977", x"7A7F8180", x"8787898D", x"8E8D8E90", x"95939190", x"93969695",
									 -- x"9A9C9B98", x"999DA09F", x"9D9D9D9F", x"A2A5A6A7", x"A7A9ACAE", x"AEAEAEAE", x"ACB0B0B1", x"B6B9BABD",
									 -- x"BDBEBFC1", x"C4C5C3BF", x"C6C7C8C8", x"C9C8C6C5", x"C9C9C9C8", x"C7C6C5C4", x"C7C8C9C8", x"C6C7C9CC",
									 -- x"CACACBCC", x"CDCDCFD1", x"D0CECED0", x"D3D5D5D4", x"D4CFD0D6", x"D6D0CED2", x"D1CDC8C7", x"C8C9C7C4",
									 -- x"C2BDBABA", x"B9B5B5B7", x"B5B3B1AF", x"AFAFACA9", x"A8A7A39E", x"9D9E9D9C", x"9A9A9490", x"918F8B8C",
									 -- x"7B7F7E7C", x"80818285", x"84878A8C", x"8D8D8D8E", x"9090908F", x"8E8D8E8E", x"908F8F91", x"92939597",
									 -- x"97989898", x"97979898", x"989A9A9A", x"9B9EA0A0", x"A09F9F9E", x"9E9FA0A1", x"A19F9E9D", x"9C9A9A9B",
									 -- x"98999999", x"97969695", x"96969797", x"94909091", x"8D8E9091", x"8F8B898A", x"8A8B8A88", x"86858687",
									 -- x"87848282", x"82807D7C", x"82828180", x"80828281", x"8383817F", x"7E7F7E7D", x"7E7B7878", x"77767778",
									 -- x"79787878", x"77777676", x"76757372", x"73767775", x"797B7A7B", x"7E7E7E82", x"8285888A", x"8D939698",
									 -- x"9A9EA09F", x"9FA2A4A3", x"A6A6A6A8", x"A9AAAAA9", x"A8A9ABB0", x"B5B8BCC0", x"C3C5C8CB", x"CECECECE",
									 -- x"D0CFCECC", x"CBCAC9C9", x"CCCCCBCA", x"C9C8C8C8", x"C8C7C5C4", x"C4C5C5C5", x"C3C4C4C4", x"C3C3C3C3",
									 -- x"C3C5C7C7", x"C7C9C9C8", x"C9CACBCC", x"CCCCCCCD", x"CFCFCECE", x"CFCFCFCE", x"CFD0D1D1", x"D1D0D0D0",
									 -- x"D0D0D1D2", x"D4D3D1CF", x"CCC9C7C5", x"C5C5C4C3", x"C5C7CACD", x"CDCED0D1", x"D3D4D6D7", x"D7D7D7D8",
									 -- x"D8D9DAD9", x"D8D8DADD", x"DCDDDFE0", x"E1E1E2E3", x"E2E4E7EA", x"EBEBEBEB", x"EEEEEEED", x"EDEFEFEF",
									 -- x"F3F3F4F5", x"F5F6F6F6", x"F4F3F2F1", x"F0EFEFEE", x"ECECECEB", x"EAE9EAEB", x"ECECECEC", x"ECECECEC",
									 -- x"ECEDEDEE", x"EEEDEBEB", x"ECEBEAE9", x"E8E7E6E6", x"E4E1E3E3", x"E0DFDEDA", x"D9D6D4D4", x"D4D2D0CF",
									 -- x"CBC7C4C2", x"C0BCB9B8", x"B5B5B3AF", x"AAA6A3A2", x"9D9B9998", x"96918A86", x"807D7C7A", x"7573726F",
									 -- x"69666362", x"62605E5B", x"5B5A5957", x"55545352", x"4E4E4F50", x"4F4E4D4C", x"4D4D4D4D", x"4B494949",
									 -- x"464A4B47", x"44454747", x"46494B4A", x"494A4C4D", x"4C4F4E4E", x"51525357", x"5556575A", x"5D5B5A5F",
									 -- x"66696C6C", x"6B6D7278", x"78797978", x"7A808382", x"88878B91", x"93929294", x"97949090", x"93989998",
									 -- x"9C9D9C99", x"999EA09F", x"9F9D9B9C", x"A1A6A8A9", x"A8A9ACAF", x"B0B1B0B0", x"B0B3B2B2", x"B6B8B9BC",
									 -- x"BEBEBDBD", x"C0C4C4C3", x"C6C8C8C7", x"C7C8C8C8", x"C8C9CAC8", x"C8C8C9C8", x"C8CACBC9", x"C7C8CACB",
									 -- x"C9C9CACC", x"CCCDD0D3", x"D1D0D0D1", x"D3D4D4D3", x"D3D4D4D3", x"D4D4D2CF", x"D1CCC6C5", x"C7C8C6C3",
									 -- x"C0BEBDBD", x"BAB6B3B1", x"B5B3B0AD", x"ACADACAA", x"A7A6A19D", x"9B9C9C9A", x"9696918F", x"908F8C8D",
									 -- x"7D7F7D7B", x"7F828284", x"8486898B", x"8B8C8C8D", x"92918E8C", x"8B8C9093", x"918F8F91", x"93939497",
									 -- x"96969695", x"94949596", x"96979798", x"9A9D9D9C", x"9D9D9E9F", x"9F9FA0A0", x"A19D9B9B", x"9C9A9999",
									 -- x"98999998", x"97959596", x"96959595", x"93909092", x"8D8D8E8E", x"8D89898A", x"8A898887", x"86868686",
									 -- x"88848283", x"84827F7E", x"7F818281", x"81828282", x"83818080", x"807E7D7D", x"7F7B7978", x"78777879",
									 -- x"79797877", x"77767675", x"75757472", x"74767674", x"797B7A7C", x"7F7E7E83", x"8384878C", x"8F929599",
									 -- x"9BA0A2A1", x"A2A5A5A3", x"A6A6A6A8", x"A9AAAAA9", x"A9AAADB1", x"B5B7BCC0", x"C4C6C9CD", x"D0D1D0CF",
									 -- x"D1D0CECC", x"CBCBCBCC", x"CDCECFCE", x"CDCBCAC9", x"CAC8C6C5", x"C5C6C6C6", x"C5C5C5C5", x"C5C5C4C3",
									 -- x"C4C6C8C7", x"C8C9CACA", x"CBCCCDCD", x"CDCDCDCD", x"D0CFCECE", x"CFCFCECD", x"D0D1D3D3", x"D3D2D2D1",
									 -- x"D1D0CFD0", x"D2D2D0CE", x"CAC8C6C6", x"C6C5C4C2", x"C6C8CBCC", x"CDCED0D2", x"D6D7D9DA", x"DADBDCDD",
									 -- x"DBDDE0DF", x"DEDDDEE0", x"DDDEE0E1", x"E2E3E4E5", x"E5E6E9EC", x"EDEDEDED", x"EEF0EFEE", x"EEF1F2F1",
									 -- x"F4F5F5F6", x"F7F7F8F8", x"F6F5F4F3", x"F2F1F0F0", x"EFEFEEED", x"EBEBECED", x"EEEDECEC", x"ECECEDEE",
									 -- x"EDEEEFF0", x"EFEEEDEB", x"EDECEAE9", x"E7E7E6E6", x"E4E1E3E4", x"E0DFDEDA", x"DCD8D5D5", x"D5D2CFCE",
									 -- x"CCC9C7C6", x"C2BDBABA", x"B7B5B2AE", x"A8A4A2A1", x"9D9B9895", x"938E8782", x"7E7A7976", x"72706F6A",
									 -- x"67656260", x"605E5B58", x"59595856", x"55535150", x"4E505152", x"514F4C4B", x"4E4C4B4C", x"4C494848",
									 -- x"44494945", x"42454746", x"4A4A4A4C", x"4C4C4C4E", x"4C505051", x"55555557", x"5858585B", x"5F5D5E65",
									 -- x"676A6E6E", x"6D6F7479", x"78787879", x"7D828586", x"8A8D8F91", x"94969796", x"95949393", x"969A9B9A",
									 -- x"9C9E9D9B", x"9CA0A19F", x"A09E9D9E", x"A1A5A7A7", x"ABABACAE", x"B0B1B0AF", x"B4B5B2B1", x"B6B7B7B9",
									 -- x"B9BBBDBD", x"BFC3C6C7", x"C3C7C9C8", x"C6C7C9C9", x"C7C9CAC9", x"C8CACBCA", x"C8CBCBC9", x"C7C9CBCC",
									 -- x"CACACCCD", x"CDCDD0D4", x"D1D2D2D3", x"D4D4D4D4", x"D4D4D4D3", x"D2D2D0CE", x"D0CCC7C6", x"C7C7C4C1",
									 -- x"BEBEBCBA", x"B8B6B3B0", x"B0B0AFAB", x"AAAAAAA8", x"A6A5A19D", x"9B9B9A98", x"9897928F", x"908F8C8D",
									 -- x"7E807C7A", x"7F828283", x"8386888A", x"8A8B8C8D", x"8D8F9091", x"90909192", x"92919193", x"94949497",
									 -- x"93939290", x"8F909192", x"96979697", x"999B9A97", x"9B9C9D9F", x"9F9E9D9C", x"A09B9798", x"9A999898",
									 -- x"97989998", x"96959697", x"94908F90", x"91909091", x"928C8787", x"8A8A8989", x"88878585", x"86878787",
									 -- x"87828081", x"82817F7E", x"7C808382", x"81828383", x"83808082", x"817D7A7B", x"7D7A7778", x"7878797B",
									 -- x"79787776", x"75757474", x"75757474", x"76787775", x"7A7B7B7C", x"7F7E7E83", x"8584888D", x"90909297",
									 -- x"9EA1A29F", x"9FA3A5A4", x"A5A5A5A6", x"A8A8A7A6", x"ABACAFB2", x"B5B7BCC0", x"C6C6C8CB", x"CED0D1D1",
									 -- x"CFCECCCB", x"CBCCCDCE", x"CCCED1D2", x"D0CECCCB", x"CAC9C7C6", x"C7C7C7C7", x"C7C6C5C5", x"C5C5C3C1",
									 -- x"C4C6C7C6", x"C7C9CAC9", x"CBCCCDCD", x"CDCDCCCD", x"CFCECECE", x"CFD0CFCE", x"D2D3D4D5", x"D4D2D1D1",
									 -- x"D2D0CFCF", x"D0D0CECD", x"C8C7C7C7", x"C7C6C3C1", x"C7C9CACB", x"CCCDD1D3", x"D6D7D8D9", x"DADBDDDE",
									 -- x"DDE0E4E4", x"E3E1E1E2", x"DFE1E2E4", x"E5E6E7E8", x"ECEDEFF0", x"F1F1F1F1", x"EEF0F0EF", x"F0F3F3F2",
									 -- x"F4F4F5F6", x"F7F7F8F8", x"F7F6F6F5", x"F3F2F2F1", x"F0F1F0EF", x"EDEDEEEF", x"EFEEECEB", x"EBECEEEF",
									 -- x"EFEFEFEE", x"EEEEEEEE", x"ECEBE9E7", x"E5E5E5E5", x"E5E2E4E4", x"E0DFDDD9", x"DBD7D4D5", x"D5D3D0CF",
									 -- x"CCCBCAC9", x"C4BEBBBA", x"B9B3ADAA", x"A9A7A29E", x"9D9B9793", x"908B8580", x"7A767473", x"70706E69",
									 -- x"6865625F", x"5E5B5855", x"56555453", x"52504D4C", x"4E4F4F4E", x"4D4B4B4A", x"4B484748", x"49464444",
									 -- x"47484643", x"454B4B46", x"4B47464B", x"4E4D4C4E", x"4C505051", x"55555355", x"5958575A", x"5E5D5F67",
									 -- x"62676D6F", x"7073787D", x"7978797D", x"8286898B", x"8D929491", x"93999A95", x"94969898", x"999C9D9C",
									 -- x"9B9E9E9D", x"9EA1A29F", x"9FA0A1A2", x"A3A3A3A2", x"AAA9A9AB", x"AFB2B2B1", x"B8B6B1B2", x"B8B9B8B9",
									 -- x"B6BCC1C1", x"C0C1C3C5", x"C0C7CDCD", x"CBCACAC9", x"C8CBCCCA", x"C9CACBCA", x"CBCECECA", x"C9CBCECF",
									 -- x"CFD0D1D2", x"D1D0D2D5", x"D1D2D4D5", x"D5D5D5D6", x"D8D1D0D5", x"D4CCCACF", x"CDCAC7C6", x"C5C3C0BE",
									 -- x"BDBDB9B3", x"B2B4B4B1", x"AAADAEAC", x"AAAAA8A5", x"A4A4A29E", x"9C9B9997", x"9B9A938E", x"8F8C898A",
									 -- x"797E7E79", x"79808382", x"83858686", x"878B8F90", x"8E8F9191", x"90919293", x"908F9093", x"96979693",
									 -- x"908F9091", x"8F8D8D90", x"8F919394", x"96989795", x"9999999B", x"9C9D9D9C", x"9E9C9894", x"95979794",
									 -- x"90919393", x"92919191", x"91919190", x"8E8E8F90", x"8E8D8A88", x"8788898A", x"89888686", x"85858585",
									 -- x"84868682", x"80818281", x"84828385", x"837F8084", x"8583807E", x"7E7D7B79", x"797A7977", x"77797979",
									 -- x"79787675", x"74737271", x"72747676", x"76767879", x"797B7E80", x"81818181", x"82838689", x"8D92979A",
									 -- x"9F9FA0A1", x"A3A5A6A7", x"A3A5A7A7", x"A8AAAAA9", x"AAB1B3B0", x"B1B8BDBC", x"C2C6CBCD", x"CECECECE",
									 -- x"D0CFCDCC", x"CDCDCCCC", x"CCD0D3D2", x"D2D2D2D0", x"CAC7C8CA", x"C8C4C3C6", x"C4C4C4C4", x"C5C5C6C6",
									 -- x"C7C7C6C4", x"C6CACAC9", x"CBCBCBCC", x"CECECDCB", x"CDCFD0D0", x"CECECFD1", x"D2D1D1D1", x"D3D4D3D2",
									 -- x"D0D1D1CE", x"CDCDCDCA", x"C9C5C6C7", x"C3C3C6C7", x"CACACACA", x"CBCDD0D2", x"D9D9DADD", x"DEDDDEE1",
									 -- x"E1E3E5E7", x"E8E7E4E2", x"E2E3E5E6", x"E7E7E8E9", x"ECEEEFEE", x"F0F2F3F2", x"F2F1F1F2", x"F3F4F4F3",
									 -- x"F6F5F5F6", x"F8F8F6F5", x"F8F6F5F5", x"F4F2F2F3", x"F3F2EFED", x"EDEEEEEE", x"EDEEEFEE", x"ECEBEDEF",
									 -- x"F0EFEEEE", x"EFEEEBE9", x"EEECE9E6", x"E5E5E6E6", x"E3E2E0DF", x"DFDEDCDB", x"D9D7D5D6", x"D5D2D0CF",
									 -- x"CEC9C9CB", x"C6C1BDB9", x"B7AFACAB", x"A6A5A4A1", x"9C9A9793", x"8D878382", x"7E7C7771", x"6E6D6A67",
									 -- x"66636360", x"5A595A57", x"56535050", x"504E4E4E", x"4D4C4C4B", x"4947484B", x"484A4A46", x"43444545",
									 -- x"49464241", x"44494947", x"47454946", x"494C464E", x"5152504F", x"50545553", x"5257595C", x"61626265",
									 -- x"6665686F", x"74777B7E", x"7B7D8185", x"888B8D8E", x"95959595", x"96989A9C", x"98989A9F", x"A09D9D9F",
									 -- x"9E9D9A9A", x"9DA1A5A8", x"9FA0A3A4", x"A19DA0A5", x"A7AAABAE", x"A8A7B2B6", x"B9B4B2B3", x"B5B4B4B7",
									 -- x"B4BAC0C0", x"BFBFC1C1", x"C4C5CACA", x"C7C7CACA", x"C9C8C7C9", x"CBCCCCCB", x"CACCCDCC", x"CACACDD1",
									 -- x"CECECECE", x"D0D2D1CF", x"D5D3CECE", x"D3D4D1D1", x"D2D0D0D0", x"D2D2CECA", x"C9C8C8C7", x"C3BEBDBE",
									 -- x"BBB9B7B5", x"B4B3B2B0", x"ACACABA8", x"A6A6A4A2", x"A0A2A19F", x"9E9D9B98", x"95959492", x"8E8B8887",
									 -- x"7A7D7C7B", x"7C818381", x"81858889", x"8A8D8E8E", x"8F909090", x"8F8F9091", x"93939395", x"97979491",
									 -- x"9391908F", x"8D8B8B8E", x"8D919493", x"92939494", x"93949698", x"98989797", x"99989491", x"93959492",
									 -- x"8F909191", x"908F8F8F", x"8C8D8F8E", x"8D8D8D8D", x"8D8C8987", x"86858687", x"87878785", x"84848688",
									 -- x"83848481", x"7F808180", x"83818285", x"84818082", x"80807F7E", x"7D7C7A79", x"7B7B7A77", x"77787978",
									 -- x"77767675", x"75757574", x"74757778", x"79797A7B", x"7A7B7B7C", x"7D7E8182", x"8284878A", x"8E929799",
									 -- x"9FA0A2A4", x"A4A5A5A6", x"A5A6A7A7", x"A8AAAAA9", x"AAAEB1B0", x"B1B7BCBE", x"C0C3C7CA", x"CBCDCED0",
									 -- x"CECCCBCB", x"CBCCCCCB", x"CED2D4D4", x"D3D3D2D1", x"CBC8C8CA", x"C9C5C5C7", x"C7C7C7C7", x"C8C8C9C9",
									 -- x"C7C8C6C4", x"C5C8CAC9", x"CACACBCC", x"CDCDCCCB", x"CCCECFCF", x"CECECFD1", x"D2D1D1D2", x"D4D4D3D3",
									 -- x"D0D1CFCD", x"CCCECECC", x"CBC7C8C9", x"C5C5C9CA", x"C9C9C9C9", x"CACCD0D3", x"D8D8D9DC", x"DEDFE2E6",
									 -- x"E6E7E8EA", x"EAE9E6E3", x"E3E4E6E7", x"E9EAECED", x"EFF0F1F1", x"F2F4F4F3", x"F4F3F3F3", x"F3F4F4F4",
									 -- x"F6F6F7F7", x"F7F6F7F7", x"F6F4F4F5", x"F5F4F4F6", x"F5F2F0EF", x"EEEEEEEE", x"EEEEEFEE", x"ECEDEFF1",
									 -- x"F2F0EFEF", x"F0EFEDEB", x"EBE9E6E4", x"E3E3E2E2", x"E1DFDDDC", x"DBDBDAD9", x"D8D7D7D7", x"D5D1CECE",
									 -- x"CBC7C8C9", x"C5C0BDB9", x"B6AFACAA", x"A5A3A2A0", x"9E9A9692", x"8B847F7E", x"7D7B7670", x"6D6B6965",
									 -- x"6460605E", x"59585855", x"524F4E4E", x"4E4D4C4C", x"4A494A4A", x"4947494B", x"45474744", x"42424241",
									 -- x"44434140", x"43474744", x"47454843", x"464B464D", x"51514F4D", x"4E515353", x"52585C5E", x"61616266",
									 -- x"6A6A6C72", x"76787A7C", x"7C7E8185", x"898D8F91", x"93959698", x"98989999", x"A0A1A2A3", x"A19E9D9E",
									 -- x"9D9EA0A1", x"A0A1A3A5", x"A5A2A1A3", x"A4A4A2A2", x"A8AAABB0", x"ADAAB1B1", x"B7B5B3B5", x"B7B8B8B9",
									 -- x"B6BCC0C0", x"BFC1C2C2", x"C3C7CACB", x"CAC9C9CA", x"CAC8C8C9", x"CBCBC9C7", x"CCCCCCCC", x"CBCCCECF",
									 -- x"CDCFD0CF", x"CFD0D0CF", x"D0D1D1D2", x"D7D5CECC", x"CFCDCCCC", x"CDCDCAC8", x"C7C5C5C5", x"C2BEBCBC",
									 -- x"BDBAB6B3", x"B2B1B1B0", x"AEACA9A7", x"A7A7A4A0", x"A3A3A09C", x"9A999693", x"9593918E", x"8C8A8989",
									 -- x"7B7A7B7D", x"81838483", x"8285898A", x"8C8E8F8E", x"8F90908F", x"8F909192", x"94939394", x"9594908D",
									 -- x"93918F8E", x"8C8A8B8E", x"8B909390", x"8D8D8F92", x"8F929596", x"95949393", x"9493908F", x"9092918E",
									 -- x"8D8D8E8D", x"8D8C8C8D", x"88898B8C", x"8C8B8B8B", x"8C8A8886", x"85858586", x"86888887", x"8586898C",
									 -- x"85848280", x"80818180", x"81808286", x"87848282", x"7E7E7E7E", x"7D7C7B7A", x"7A7A7976", x"75777877",
									 -- x"77777777", x"78787777", x"7878797B", x"7D7D7D7C", x"7C7C7C7C", x"7D7F8284", x"8385888C", x"8F929698",
									 -- x"9EA1A4A6", x"A5A4A4A5", x"A7A8A8A7", x"A7AAABAA", x"ABADAFB0", x"B1B5BABE", x"BFC1C4C6", x"C8CACDCF",
									 -- x"CCCBCACA", x"CBCCCCCC", x"CDD0D2D3", x"D3D2D1D0", x"CFCBCACB", x"CBC8C8CA", x"C9C9C9C9", x"C9C9C9C9",
									 -- x"C8C8C7C5", x"C4C6C8C9", x"C9CACBCB", x"CBCBCCCC", x"CBCDCECF", x"CECFD0D2", x"D2D2D2D3", x"D4D4D3D2",
									 -- x"D1D0CECC", x"CDCFCFCD", x"CAC6C7C9", x"C6C6CACA", x"C9C9C9C8", x"C9CCD1D5", x"D7D8DADE", x"E0E2E5E8",
									 -- x"E9E9E9EB", x"ECEBE7E4", x"E4E5E6E7", x"E9ECEDEF", x"F0F2F3F2", x"F3F5F5F4", x"F6F5F3F3", x"F3F4F4F3",
									 -- x"F5F6F7F6", x"F4F4F6F8", x"F5F4F5F6", x"F7F6F6F7", x"F6F3F0F1", x"F0EDEDEF", x"EEEEEFEE", x"EDEEF0F2",
									 -- x"F2F0EEEE", x"EEEDEBE9", x"E8E6E4E3", x"E2E1E0DF", x"DFDDDBDA", x"D9D9D8D8", x"D6D6D7D7", x"D4CFCBCB",
									 -- x"C8C4C5C7", x"C3C0BDB8", x"B5AEABA9", x"A4A1A09D", x"9E99948F", x"8A847F7D", x"7C79746E", x"6B696663",
									 -- x"635F5E5D", x"5A595955", x"504E4D4E", x"4E4B4A4A", x"4A494949", x"46444446", x"45464544", x"4343413F",
									 -- x"40404040", x"42444442", x"46474742", x"454B484C", x"51525250", x"50525354", x"545B5F61", x"62626469",
									 -- x"70707276", x"797A7C7E", x"7F828588", x"8B8E9192", x"94969899", x"9999999A", x"9FA3A4A2", x"A09FA0A1",
									 -- x"9CA1A5A6", x"A3A1A3A5", x"A8A5A3A3", x"A6A8A5A1", x"AAAAA9AF", x"AEACB0AC", x"B0B0B1B2", x"B5B8B9B7",
									 -- x"B9BCBEBF", x"C0C2C2C2", x"C4C9C7C8", x"CDCBC8CC", x"CBC9C8CA", x"CCCCC9C5", x"CCCCCBCB", x"CBCCCCCC",
									 -- x"C9CDD0D0", x"CECFCFCF", x"D0D1D0D0", x"D3D2CECF", x"D0CECDCC", x"CBCAC8C7", x"C4C2C2C2", x"C1BEBBB9",
									 -- x"BEBAB5B1", x"AFAFAFAF", x"ACA9A6A4", x"A6A7A39E", x"A09E9A96", x"96979593", x"92908D8B", x"8B8A8988",
									 -- x"7C797A7F", x"83848588", x"85878989", x"8B8E9090", x"8F8F9090", x"91939495", x"94939292", x"93928F8D",
									 -- x"91908E8D", x"8C8C8D8E", x"898D8F8D", x"89898C8F", x"8E909393", x"91909091", x"92908F8E", x"8F8F8D8B",
									 -- x"8A8A8A8A", x"89898A8A", x"8688898A", x"8A8A8989", x"8A898786", x"86868788", x"86878787", x"8687898B",
									 -- x"87858382", x"82838281", x"80808387", x"88868586", x"81807E7E", x"7E7E7C7A", x"7B7B7976", x"76787979",
									 -- x"7B7A7A7A", x"7A7A7978", x"7B7B7C7E", x"80807F7E", x"7D7E7F80", x"80818283", x"84868A8D", x"90929596",
									 -- x"9B9FA4A5", x"A4A3A4A5", x"A8A9A8A7", x"A7AAACAC", x"AFADAEB1", x"B2B3B7BD", x"BFC0C2C4", x"C5C6C8CB",
									 -- x"CCCCCBCC", x"CCCDCDCE", x"CACCCFD1", x"D1D1D0CF", x"D0CCCACB", x"CBCACACB", x"CBCBCACA", x"C9C8C8C7",
									 -- x"C9C9C9C6", x"C5C6C8CA", x"C9CACBCB", x"CBCACBCD", x"CCCDCECF", x"CFD0D1D2", x"D3D3D3D4", x"D4D3D2D1",
									 -- x"D1D0CECD", x"CECFCECD", x"CAC6C7C9", x"C7C7CACA", x"C9CACBCA", x"CACDD2D6", x"D8DADEE2", x"E4E4E5E6",
									 -- x"E9E8E8EA", x"ECECE9E5", x"E5E5E5E6", x"E8EAECED", x"F0F2F3F2", x"F3F5F5F3", x"F6F5F3F2", x"F3F3F4F4",
									 -- x"F4F5F4F3", x"F3F3F5F6", x"F6F6F6F7", x"F6F5F5F5", x"F6F2F0F2", x"F1EEEDF0", x"EEEEEEED", x"ECEDEFF1",
									 -- x"F1F0EEEC", x"EBEAE8E7", x"E6E6E4E4", x"E3E1E0DE", x"DEDCDBDA", x"DAD9D8D7", x"D4D4D4D4", x"D1CBC9C8",
									 -- x"C5C2C3C4", x"C1BFBDB8", x"B4AEABA9", x"A39F9E9C", x"9B96908D", x"8A85817F", x"7B78736D", x"6A686562",
									 -- x"615D5B5B", x"59595853", x"504F4F4F", x"4E4A4847", x"49484747", x"44414143", x"46454343", x"4343413F",
									 -- x"3F40403F", x"40424341", x"44484844", x"474C4C4D", x"4D505253", x"53525353", x"585E6162", x"6566686E",
									 -- x"7274777A", x"7D7E8082", x"84868A8C", x"8E8F9192", x"98989899", x"999A9C9E", x"9DA2A4A1", x"9EA0A2A2",
									 -- x"9EA2A5A6", x"A4A3A5A7", x"A4A6A6A3", x"A4A7A8A5", x"ABA9A7AC", x"ABAAB0AC", x"B2B4B4B4", x"B8BDBEBB",
									 -- x"B9BABCBE", x"C0C1C1C0", x"C7C9C1C1", x"CCCDC9CF", x"CBC9C9CB", x"CFCFCBC7", x"CDCDCDCD", x"CCCBCBCB",
									 -- x"C7CACECE", x"CFCFCFCE", x"D0D1CECD", x"CFCFCED1", x"D0CFCECD", x"CBC8C7C7", x"C3C1C0C0", x"C1BFBAB7",
									 -- x"BAB8B5B2", x"AFADADAC", x"A7A5A2A1", x"A3A4A19D", x"9C999594", x"94959492", x"8D8C8B8B", x"8C8A8683",
									 -- x"7C7A7C80", x"81808489", x"8688898A", x"8C8F9190", x"90909091", x"93949696", x"94939292", x"93939392",
									 -- x"90908F8E", x"8E8E8D8C", x"888A8B89", x"88898B8B", x"8C8D8F8E", x"8C8C8D8F", x"92908F8F", x"8F8D8B8A",
									 -- x"89898A89", x"88888989", x"88888888", x"88888888", x"88878685", x"85868788", x"86858585", x"87878786",
									 -- x"89868383", x"83838383", x"80828587", x"86858687", x"86827D7C", x"7E7E7C78", x"7B7C7B79", x"797C7D7D",
									 -- x"7D7C7C7C", x"7C7C7B7B", x"7F7E7E80", x"82828180", x"7F808081", x"81828384", x"86888B8E", x"91939596",
									 -- x"999DA1A2", x"A2A2A4A7", x"A8A9A8A7", x"A8ABADAD", x"B0AEAEB2", x"B3B3B6BC", x"BEBEC1C3", x"C4C3C5C8",
									 -- x"CBCBCCCD", x"CDCDCDCD", x"CBCCCED0", x"D0D0CECE", x"CECCCACA", x"CAC9CACB", x"CCCCCCCC", x"CBCBCAC9",
									 -- x"CBCACAC8", x"C7C6C9CB", x"C9CACCCC", x"CBCBCCCD", x"CECECFD0", x"D0D1D2D2", x"D3D4D4D3", x"D3D2D1D1",
									 -- x"D2D0CFD0", x"D0CFCDCB", x"CCC8C9CB", x"C9CACCCC", x"CACBCDCD", x"CDCFD3D6", x"DBDDE0E2", x"E3E5E6E6",
									 -- x"E8E8E8E9", x"EBEBE9E6", x"E6E4E3E4", x"E6E9ECED", x"F0F2F3F3", x"F4F5F5F3", x"F6F5F3F3", x"F3F4F5F5",
									 -- x"F6F4F2F2", x"F3F4F4F4", x"F5F6F6F5", x"F5F4F3F2", x"F3F0EFF1", x"F1EFEEF0", x"EEEEEDEC", x"EBEBECED",
									 -- x"F0EFEDEC", x"EBEAE9E8", x"E5E5E4E4", x"E3E2DFDE", x"DCDCDCDC", x"DBDAD7D6", x"D4D2D1D0", x"CECAC8C8",
									 -- x"C3C1C2C2", x"BFBEBDB7", x"B3ADAAA8", x"A29E9D9A", x"97928D8B", x"89858180", x"7A78736D", x"6A686562",
									 -- x"5E5A5959", x"56565550", x"4F4E4E4F", x"4D494747", x"44434344", x"42414245", x"44413E3E", x"40403F3D",
									 -- x"3F403F3D", x"3E414241", x"42484746", x"4A4D4D4D", x"4A4B4D4F", x"4F4F5153", x"5B5F5F60", x"66696B71",
									 -- x"7375797B", x"7E808283", x"86898D90", x"91919292", x"97979899", x"9A9B9D9F", x"A1A6A7A2", x"9E9EA0A0",
									 -- x"A1A2A4A6", x"A7A6A5A5", x"A2A4A3A1", x"A3A7A9A7", x"A8A8A7AD", x"ABA9B0AE", x"B3B4B4B3", x"B7BCBEBB",
									 -- x"B9BABCBF", x"C1C1C0BF", x"C6C6BDBE", x"CCCDC8CE", x"CAC9C9CB", x"CECFCBC8", x"CCCECFCF", x"CDCCCED0",
									 -- x"C9CBCDCE", x"D0D1D0CD", x"CDD0CFCE", x"D0CDC9CA", x"CAC9CACB", x"CAC6C4C4", x"C2C0BFBF", x"C0BEB9B5",
									 -- x"B5B5B4B3", x"B0ADAAA9", x"A4A4A2A0", x"9F9F9D9B", x"9D9A9694", x"93918E8C", x"8C8A898A", x"8A878380",
									 -- x"7E7D7E80", x"7F7E8186", x"85888A8C", x"8E91908E", x"90909192", x"94959595", x"94939292", x"93949494",
									 -- x"91929291", x"908F8C89", x"88898887", x"888A8B89", x"8C8D8D8C", x"8B8B8D8E", x"918F8E8F", x"8E8C8A89",
									 -- x"89898A8A", x"89888989", x"89888686", x"86878787", x"86858483", x"83838485", x"89878586", x"89898886",
									 -- x"88858382", x"82818283", x"83848485", x"85848484", x"87837E7C", x"7D7E7B79", x"797A7A79", x"7A7D7E7E",
									 -- x"7E7D7D7D", x"7E7F8080", x"82828283", x"84848484", x"86858483", x"8385878A", x"898B8E91", x"93959798",
									 -- x"9A9C9FA1", x"A1A2A4A7", x"A7A9A9A8", x"A9ABADAC", x"AFADAEB2", x"B3B4B7BB", x"BBBBBEC2", x"C2C1C2C6",
									 -- x"C7C9CBCC", x"CCCCCBCB", x"CCCBCBCD", x"CDCCCACA", x"CDCECECD", x"CCCCCCCD", x"CBCBCCCC", x"CCCCCCCB",
									 -- x"CCCACAC9", x"C9C8C9CB", x"C9CACBCC", x"CCCCCBCB", x"CFCFD0D0", x"D1D2D2D2", x"D2D2D2D2", x"D1D0D1D1",
									 -- x"D2D1D1D2", x"D0CDCBCB", x"CBC7C8CA", x"C9C9CBCA", x"CBCBCCCD", x"CFD1D5D7", x"DDDEDFDF", x"E0E4E7E8",
									 -- x"E9E9E9EA", x"EAE9E8E7", x"E6E4E2E3", x"E6EAEDEE", x"EFF1F3F3", x"F4F6F6F4", x"F5F4F3F4", x"F5F6F6F6",
									 -- x"F6F4F2F1", x"F3F4F4F3", x"F2F3F3F2", x"F2F2F2F0", x"EFEEEEEF", x"F0F0EFEE", x"EDEDECEB", x"EAEAE9E9",
									 -- x"EAEAEAE9", x"E9E8E8E8", x"E4E3E3E2", x"E2E0DEDC", x"DADBDCDC", x"DCDAD7D4", x"D5D2CFCD", x"CCC9C7C7",
									 -- x"C2C0C0C0", x"BDBDBBB5", x"B0ABA9A7", x"A09C9B99", x"94908C8A", x"86827E7D", x"7A77726D", x"6A686662",
									 -- x"5F5B5A5A", x"56555450", x"4C4C4C4C", x"4B484849", x"45444343", x"41404144", x"423F3C3D", x"3E3F3E3E",
									 -- x"3F3E3C3B", x"3D404140", x"42474548", x"4C4B4D4D", x"4D4B4B4C", x"4D4F5357", x"5C5F5E60", x"666A6D72",
									 -- x"73767A7C", x"7D808282", x"868A8E91", x"92929495", x"9396999B", x"9C9C9C9D", x"A1A4A4A1", x"9E9E9FA0",
									 -- x"A3A3A4A7", x"AAA9A5A0", x"A5A29E9F", x"A5AAA9A5", x"A5A8AAB0", x"AEABB1AF", x"B1B0B0B0", x"B3B7B8B7",
									 -- x"BBBBBCBF", x"C1C0C0C0", x"C2C1BEC2", x"CBCAC6C9", x"C9C8C8C9", x"CBCCCAC8", x"C8CBCDCD", x"CBCBCED1",
									 -- x"CECECDCD", x"CFD0CECB", x"CFD1CDCA", x"CBC9C6C8", x"C6C5C5C8", x"C9C5C3C3", x"C0BFBDBC", x"BDBCB8B3",
									 -- x"B0B1B2B2", x"AFABA8A6", x"A4A5A39F", x"9D9C9A98", x"9A979594", x"928E8C8B", x"8C8A8785", x"8483807F",
									 -- x"7F808081", x"82828385", x"86888A8B", x"8E91918E", x"91919294", x"96979695", x"95959595", x"94949392",
									 -- x"94959492", x"91908C88", x"88898887", x"888A8A89", x"8B8B8B8B", x"8C8C8D8D", x"8D8B8B8D", x"8C8A898A",
									 -- x"87888988", x"88878787", x"87868484", x"84858585", x"83838282", x"82828383", x"8A888686", x"88898988",
									 -- x"87848282", x"817F8083", x"86858384", x"87888582", x"8583807F", x"7E7E7D7C", x"787A7B7A", x"7C7E7F7E",
									 -- x"82818081", x"82848586", x"84858686", x"8788898A", x"8A8A8988", x"87898B8D", x"8C8E9193", x"9597999B",
									 -- x"9D9EA0A2", x"A2A3A4A5", x"A7A9A9A9", x"AAABACAB", x"ADADAFB1", x"B3B4B6B8", x"B9B8BBBF", x"C0BEC0C4",
									 -- x"C4C7CACC", x"CCCBCACA", x"CBC8C8C9", x"CAC9C9CA", x"CDCFD1D1", x"CFCDCECE", x"CCCCCDCE", x"CECDCCCC",
									 -- x"CCC9C9CA", x"CAC9C9CA", x"C8C9CACC", x"CDCCCBC9", x"CECECFD0", x"D1D2D3D3", x"D0D0D0D0", x"CFCFD1D2",
									 -- x"D2D2D2D2", x"CFCCCBCD", x"CAC6C6C9", x"C8C8C9C8", x"CAC9C9CA", x"CED2D6D7", x"DBDDDEDE", x"DFE2E4E4",
									 -- x"E7E8E9E9", x"E8E8E8E8", x"E6E4E1E2", x"E5E9ECED", x"EDF0F2F2", x"F3F5F5F3", x"F3F3F2F3", x"F4F5F5F5",
									 -- x"F4F3F1F1", x"F1F2F2F2", x"F0F1F1EF", x"EEF0F0EE", x"EBEEEEEC", x"EDF0EFEB", x"ECECEBEA", x"EAE9E8E7",
									 -- x"E6E7E7E7", x"E6E5E5E4", x"E2E2E1E1", x"E0DFDDDB", x"DBDBDCDC", x"DCDAD7D5", x"D5D0CBCA", x"C9C7C4C3",
									 -- x"C1BFBFBE", x"BBBBB9B3", x"AEA9A7A5", x"9E9A9997", x"93908D8A", x"857F7C7B", x"7977726D", x"6A696663",
									 -- x"615E5E5D", x"57555451", x"4C4B4A4B", x"4947484A", x"4A484644", x"413F4043", x"413F3E3F", x"41404041",
									 -- x"3F3D3B3B", x"3E424341", x"4549444A", x"4E494D4F", x"52504E50", x"5354575B", x"5C606163", x"686A6D73",
									 -- x"73787C7D", x"7F818484", x"888B8F91", x"91929597", x"95979A9D", x"9D9D9D9D", x"A0A0A1A2", x"A1A0A1A3",
									 -- x"A6A5A5A7", x"AAAAA6A2", x"A8A29FA0", x"A5A7A7A6", x"A6A8A9B0", x"AEACB2AF", x"B4B2B2B4", x"B7B8B8B9",
									 -- x"BCBBBBBE", x"BFBEBFC1", x"C0C0C2C6", x"C6C3C4C8", x"C7C7C7C8", x"C9CBCCCC", x"CACBCCCB", x"CACACCCE",
									 -- x"CECECDCB", x"CBCCCBCA", x"CFCFC9C6", x"C8C8C7CA", x"C8C4C3C6", x"C7C3C0C0", x"BCBCBBB9", x"B9B9B6B2",
									 -- x"ADAFAFAE", x"ABA8A5A4", x"A4A3A09D", x"9C9B9895", x"93929292", x"8F8C8C8D", x"88888684", x"817F7D7C",
									 -- x"80818283", x"86888886", x"89898989", x"8C909291", x"90919295", x"98999998", x"99999999", x"98969392",
									 -- x"95969492", x"91908D89", x"888A8A89", x"888A8A89", x"87878889", x"8A8B8A89", x"8987888A", x"8B89898A",
									 -- x"84858687", x"86858484", x"85848282", x"83848483", x"81818181", x"82838484", x"87868483", x"83848789",
									 -- x"87848382", x"807F8084", x"88858285", x"8B8D8882", x"83848482", x"807F7F80", x"7B7D7E7E", x"7F828281",
									 -- x"86858484", x"8688898A", x"86878889", x"898A8D8F", x"88898A8B", x"8B8B8B8B", x"8E909295", x"97999C9D",
									 -- x"A0A1A2A4", x"A4A4A4A3", x"A7A9AAAA", x"AAABABA9", x"ADAFB0B0", x"B1B4B5B4", x"B9B7B9BD", x"BEBCBEC3",
									 -- x"C2C5CACD", x"CDCCCBCB", x"CAC8C7C9", x"CBCBCCCD", x"C9CDD1D0", x"CDCBCCCD", x"D1D1D1D1", x"D0CFCECD",
									 -- x"CBC8C7CA", x"CBC9C8C9", x"C8C8C9CB", x"CDCDCAC8", x"CDCDCECF", x"D1D3D3D3", x"CECECECE", x"CECFD2D4",
									 -- x"D2D2D3D2", x"CECACBCF", x"CBC7C7CA", x"C9C9CAC8", x"C9C7C5C8", x"CDD3D6D8", x"D7DCDFE0", x"E1E1E0DE",
									 -- x"E4E6E8E8", x"E7E7E8EA", x"E8E4E1E0", x"E3E7EAEB", x"EBEDF0F0", x"F2F4F3F2", x"F1F1F1F1", x"F2F3F2F2",
									 -- x"F0F1F1F0", x"EEEEEFF1", x"F0F1F0ED", x"ECEDEDEC", x"E9EDEEEB", x"EBF0EFE9", x"EBEBEAEA", x"EAE9E7E6",
									 -- x"E8E8E9E8", x"E6E5E3E3", x"E2E1E1E0", x"E0DEDDDB", x"DDDDDDDD", x"DCDBD9D7", x"D3CEC9C8", x"C7C4C1BE",
									 -- x"C0BEBEBD", x"B9B9B7B1", x"ACA7A6A4", x"9C989795", x"92908E8B", x"857F7C7B", x"7876716C", x"6A696663",
									 -- x"615E5F5D", x"57545350", x"4D4C4B4A", x"4847484A", x"49484645", x"42414347", x"403E3E41", x"42404041",
									 -- x"3F3D3B3C", x"41454643", x"494B444C", x"50484D51", x"54525256", x"5959595A", x"5C636667", x"6A6B6E75",
									 -- x"74797E7F", x"81848787", x"8A8D9090", x"90919498", x"9A9A9C9C", x"9D9E9FA0", x"A4A2A3A6", x"A5A3A3A6",
									 -- x"A8A5A4A5", x"A7AAAAA9", x"A8A5A4A4", x"A3A2A4AA", x"A9A8A7AC", x"ABABB2B0", x"B2AFB0B4", x"B7B5B5B6",
									 -- x"BCBABABB", x"BBBBBEC2", x"C0C0C5C7", x"C1BEC3CA", x"C6C6C7C8", x"C9CCCED1", x"D1D0CECD", x"CCCCCDCD",
									 -- x"CACCCBC8", x"C6C7C9CA", x"C7C9C8C9", x"CCCBC7C7", x"CBC5C1C4", x"C4C0BCBC", x"B8B9B8B6", x"B6B7B5B2",
									 -- x"ADAEADAB", x"A7A5A3A3", x"A19F9C9A", x"9B9C9893", x"91909090", x"8C898A8D", x"84858684", x"817D7A78",
									 -- x"81808083", x"8484878A", x"88888889", x"8B8D8F91", x"8E8C9399", x"96989D9C", x"9A9B9A98", x"96959697",
									 -- x"96969695", x"93918E8D", x"898A8A8B", x"8B8B8A89", x"8987888A", x"8A888687", x"85848587", x"86838182",
									 -- x"83838180", x"81848584", x"80828080", x"83828082", x"817F7D7E", x"7D7E8287", x"83858686", x"85858789",
									 -- x"88868484", x"83828486", x"84868788", x"8B8B8680", x"84858584", x"82818181", x"7D7D7D7F", x"83858787",
									 -- x"8784878A", x"88898E8F", x"8E8B8A8A", x"8D8F9090", x"8D8E8E8F", x"8F8F8E8D", x"8F909396", x"999CA0A2",
									 -- x"A2A4A4A3", x"A4A6A7A6", x"A7A8AAAB", x"ABABACAC", x"B0AEAEB0", x"B1B2B4B7", x"B6B6B8BB", x"BDBDC0C3",
									 -- x"C2C4C7CA", x"CCCBCAC9", x"CAC9C8C9", x"CACCCCCC", x"CDCDCDCD", x"CCCDCECF", x"CFD2D4D3", x"D2D1CFCC",
									 -- x"CCCAC8C7", x"C8CACBCB", x"C8C9CACB", x"CCCBCBCA", x"CBCED1D1", x"D0D0D0D1", x"CDCCCCCD", x"CECED2D5",
									 -- x"D3D2D2D3", x"D1CDCBCB", x"CCC8C8C9", x"C4C3C6C7", x"C6C6C7C7", x"C8CBD0D5", x"D3D5D6D6", x"D7DADBDA",
									 -- x"DBDEE2E5", x"E7E7E8E9", x"E9E7E3E0", x"E0E3E7EA", x"E9EBEFF0", x"F0F0F1F2", x"F3EFEBED", x"EFEFEFEF",
									 -- x"F3EFEBEB", x"EDEFEFED", x"F0F1F1EF", x"ECEAEBEC", x"EEEDEAE9", x"E8E9EAEB", x"EEEAE9EA", x"EAE7E8EC",
									 -- x"E5E5E4E4", x"E4E4E3E3", x"E1E3E2DE", x"DDDEDEDD", x"DEDDDCDB", x"DBDAD9D8", x"D1CCC6C3", x"C2C1BEBC",
									 -- x"BDBCBAB9", x"BBBBB5AF", x"AAA8A5A0", x"9C999797", x"8F8B8887", x"86827E7D", x"79746F6D", x"6B666363",
									 -- x"5F5E5D5A", x"56535150", x"4E4A4849", x"48454649", x"4A464241", x"43454442", x"3F3F4041", x"42403C3A",
									 -- x"3A3C393A", x"42474543", x"49494A4C", x"4E4F4E4D", x"51535556", x"585C5D5D", x"5E646869", x"6B6F7374",
									 -- x"747A7E80", x"81818690", x"8A8E9395", x"9596999C", x"9D9F9D99", x"999FA3A3", x"A5A1A0A3", x"A4A3A4A8",
									 -- x"A3A4A5A7", x"A6A5A6A8", x"A3A6A8A7", x"A4A5ABB1", x"A8A8A7AA", x"B0B2B2B6", x"AFAFB2B5", x"B5BABBB6",
									 -- x"B8BCC0BF", x"BDBDBEBE", x"BEC2C5C5", x"C2C1C4C7", x"C6C7C8C8", x"C8CACDCF", x"CBCACBCC", x"CBC9C9CA",
									 -- x"CBC9C9C9", x"C8C5C5C5", x"C6C6C6C7", x"C8C9C8C7", x"C0C2C2BE", x"BDBFBDB8", x"B7B4B7BB", x"B7B2B0AF",
									 -- x"B2ADAAAA", x"A8A3A09F", x"A09E9C99", x"97969392", x"918E8E90", x"8D888688", x"8185837D", x"797A7A79",
									 -- x"84838384", x"84838487", x"8A898888", x"898A8C8E", x"9090959A", x"9A9A9D9E", x"9D9C9B9A", x"98979797",
									 -- x"95959595", x"9593918F", x"8B8A8A8A", x"8C8C8A88", x"87858586", x"87868687", x"88868587", x"8783807F",
									 -- x"7F81817F", x"7D7F8080", x"82848280", x"82807C7D", x"7A79797B", x"7C7D8185", x"84868787", x"8787888A",
									 -- x"87878787", x"84828487", x"85868686", x"898A8783", x"85858584", x"83838282", x"81808183", x"8688898A",
									 -- x"89878A8D", x"8B8C9090", x"95939190", x"92939292", x"91919091", x"91929191", x"91939597", x"9A9DA0A2",
									 -- x"A2A4A5A5", x"A6A8A9A8", x"A8A9AAAB", x"ACACADAE", x"ACACAEB2", x"B4B4B5B6", x"B6B7B8BB", x"BBBBBDC0",
									 -- x"C1C2C4C6", x"C8C8C8C8", x"C8C7C7C8", x"CACBCCCC", x"CCCCCDCC", x"CCCDCFD0", x"D1D4D5D4", x"D3D1CFCD",
									 -- x"CCCAC8C7", x"C8C9C9C9", x"C8C9CACB", x"CBCCCBCB", x"CBCDCFCF", x"CECDCECF", x"CECDCDCE", x"CDCDCFD2",
									 -- x"D2D2D4D4", x"D1CCCBCC", x"CCC7C8C8", x"C4C3C6C6", x"C0C1C1C1", x"C2C5C9CC", x"D0D2D4D5", x"D7DADBDA",
									 -- x"D7DBE0E3", x"E5E5E6E7", x"E7E5E2E0", x"E0E2E5E7", x"E8EAEDEE", x"EEEEEFF0", x"F0ECEAEB", x"ECEBEAEB",
									 -- x"EFECEAE9", x"EBEDEDEC", x"EDEFF0EF", x"EDECEDEE", x"ECECEBEA", x"EAEAEBEC", x"EEEBEAEB", x"EAE7E7E9",
									 -- x"E8E7E6E6", x"E5E4E3E2", x"E1E2E1DF", x"DEDFE0DF", x"DCDCDCDC", x"DBD9D6D4", x"D2CEC9C3", x"BFBCBAB9",
									 -- x"B8BAB9B8", x"B7B6B3B0", x"AAA7A39F", x"9C999694", x"8F8A8786", x"85807B78", x"76726F6D", x"6A656261",
									 -- x"5E5B5856", x"5553504E", x"4E4C4A4A", x"49474748", x"48454241", x"43454544", x"43424041", x"42403C38",
									 -- x"3A40403E", x"40414245", x"49494A4D", x"4F4F4E4D", x"55565859", x"5A5B5D5F", x"5E626668", x"6A6E7172",
									 -- x"7879797C", x"8386888D", x"8D8F9191", x"9193979C", x"9A9C9C98", x"999EA1A1", x"A3A0A0A3", x"A4A2A3A5",
									 -- x"A7A7A9AB", x"A9A6A6A7", x"A5A7A7A5", x"A2A3A8AD", x"ACAEAEAE", x"B0AEAEB3", x"B7B5B5B5", x"B4B8BCB9",
									 -- x"B9BCBFBE", x"BDBEC0C0", x"BDC0C4C4", x"C2C2C5C8", x"CBCAC8C7", x"C7C7C8C8", x"CBCACACA", x"C8C6C6C8",
									 -- x"C9C7C5C6", x"C6C5C4C4", x"C3C3C4C4", x"C3C3C4C5", x"BEBEBEBF", x"BDBAB7B5", x"B8B3B4B7", x"B3AFB0B0",
									 -- x"ADAAA6A5", x"A4A2A09E", x"9D9C9B98", x"95939291", x"908C8B8C", x"89848284", x"827F7B77", x"75747576",
									 -- x"83828385", x"8686888A", x"8A898887", x"87898B8C", x"8F93969A", x"9D9C9CA0", x"9E9D9C9B", x"9A999897",
									 -- x"99989696", x"9694908D", x"8D8B8989", x"8A898785", x"87848383", x"84848485", x"86848385", x"87858280",
									 -- x"7C7F807D", x"7A797A7B", x"8183817F", x"7F7C7879", x"7575777A", x"7C7E8184", x"85858687", x"88888888",
									 -- x"87888A8A", x"86838588", x"87868585", x"87898986", x"88878685", x"86868685", x"85858587", x"898B8C8C",
									 -- x"8D8B8F93", x"91919495", x"97959495", x"96979796", x"96959494", x"94959595", x"9597989A", x"9C9FA1A3",
									 -- x"A4A6A8A8", x"A9ABABAA", x"AAAAABAC", x"ADAEAFAF", x"ABABADB1", x"B3B3B3B5", x"B5B6B7BA", x"BABABBBD",
									 -- x"BFC0C1C2", x"C3C4C5C6", x"C6C6C6C7", x"C9CBCCCC", x"CBCBCCCC", x"CDCDCFD1", x"D2D4D5D3", x"D1D0CECC",
									 -- x"CCCBC9C9", x"C8C8C8C8", x"C8C9C9CA", x"CBCCCCCC", x"CBCDCDCD", x"CCCBCCCD", x"CDCCCDCE", x"CDCCCCCE",
									 -- x"CFD1D4D4", x"CFCBCBCD", x"CBC6C6C7", x"C4C5C6C5", x"C3C3C3C4", x"C5C7C9CA", x"CCCED1D3", x"D6D9DAD9",
									 -- x"D6DADFE4", x"E5E6E6E6", x"E4E3E1E0", x"E0E1E3E4", x"E6E8EAEB", x"EBEBECEC", x"ECEAE9E9", x"E8E7E6E7",
									 -- x"EBEBEAEA", x"EAEAEBEB", x"EBEDF0F0", x"EFEEEEEE", x"ECECECEC", x"ECECECEC", x"EEECEBEC", x"EBE7E6E8",
									 -- x"E9E9E8E7", x"E6E5E4E3", x"E0E1E1DF", x"DEDFE0E0", x"DDDEDEDF", x"DDD9D5D2", x"D0CDC9C4", x"BFBCBCBC",
									 -- x"B7BABAB8", x"B4B2B1B0", x"AAA6A19D", x"9A979390", x"8D898584", x"837F7975", x"7573706E", x"6A666463",
									 -- x"5F5C5856", x"5654514F", x"4C4C4B4A", x"4A4A4948", x"46444343", x"43454646", x"48454141", x"42413D38",
									 -- x"3F403E3D", x"43454343", x"47484A4E", x"51525251", x"5555585B", x"5B595C60", x"60636668", x"6C707273",
									 -- x"7A7A797D", x"8588898E", x"90909190", x"9093979B", x"9A9D9D9B", x"9CA0A2A2", x"A19F9FA2", x"A3A1A0A2",
									 -- x"A2A4A7AA", x"A9A6A5A6", x"A6A7A6A5", x"A3A4A8AB", x"A9AEB0B1", x"B1ADAEB4", x"B8B6B7B6", x"B3B7BAB9",
									 -- x"BBBCBDBD", x"BEC0C2C2", x"C0C3C5C4", x"C2C1C2C4", x"CAC8C7C7", x"C9C9C8C7", x"CAC9C8C7", x"C6C4C5C7",
									 -- x"C7C4C2C3", x"C4C3C3C3", x"C0C1C2C1", x"BFBEC0C2", x"BFBCBCBF", x"BDB6B4B7", x"BAB5B5B7", x"B2AFAFAE",
									 -- x"A8A6A3A0", x"A0A09F9D", x"999A9996", x"928F8F90", x"8D8A8888", x"85807E7F", x"827A7676", x"76727274",
									 -- x"83828386", x"89898A8C", x"8A898888", x"88898B8B", x"8B929497", x"9E9D9CA2", x"A09F9E9E", x"9F9E9C9A",
									 -- x"9D9A9897", x"9795908C", x"8F8E8C8A", x"89888686", x"88868483", x"83828282", x"83828384", x"85848280",
									 -- x"7C7E7E7B", x"78787878", x"7B7E7D7B", x"7C797677", x"7676787A", x"7D7F8183", x"84848586", x"88888887",
									 -- x"89898A8A", x"87858688", x"88878686", x"888A8988", x"8B898887", x"88888888", x"8888898A", x"8B8C8C8C",
									 -- x"908F9397", x"95969A9B", x"9999999A", x"9B9B9B9A", x"9C9B9999", x"99999999", x"989A9C9E", x"A0A2A4A6",
									 -- x"A8AAABAB", x"ACADACAA", x"ACABABAC", x"ADAEAFAF", x"B0AEAEAF", x"B0B1B3B5", x"B4B4B6B9", x"BABABBBD",
									 -- x"BEBEBFC0", x"C1C2C4C4", x"C6C6C7C8", x"C9CACBCB", x"CBCBCBCD", x"CDCDCFD1", x"D0D2D3D1", x"CFCECCCA",
									 -- x"CCCBCACA", x"C9C8C8C8", x"C8C8C9C9", x"CACCCCCD", x"CCCDCDCC", x"CBCACBCC", x"CCCCCCCE", x"CECCCCCD",
									 -- x"CDCFD1D1", x"CECCCBCC", x"CAC5C5C6", x"C4C5C6C3", x"C1C1C1C3", x"C4C5C6C5", x"C8CBCFD1", x"D4D7D8D7",
									 -- x"D5D9DFE3", x"E4E4E4E4", x"E2E1E0DF", x"DFE0E1E3", x"E3E5E8EA", x"E9E9E9E9", x"EAEAEAE9", x"E7E6E6E7",
									 -- x"EAECECEB", x"EAE9EAEB", x"EBEDEFF1", x"F0EFEDED", x"EEEEEDED", x"ECECECEC", x"EFEDECEC", x"EBE8E7E9",
									 -- x"E8E8E7E7", x"E7E6E4E3", x"E0E1E1DF", x"DEDEDFDF", x"DFDFDFDF", x"DDD9D4D0", x"CDCAC6C1", x"BEBCBBBB",
									 -- x"B8B9B8B5", x"B1AEADAD", x"A9A59F9B", x"9995918D", x"8C878382", x"817F7A75", x"7674716D", x"6A666565",
									 -- x"605E5A58", x"56545251", x"4B4C4B48", x"494C4C48", x"45454545", x"44454647", x"49464342", x"43423F3C",
									 -- x"3E3E3B3E", x"474A4847", x"484A4C4F", x"52535455", x"5453575C", x"5B595C63", x"62636669", x"6E727475",
									 -- x"777B7D80", x"8485888F", x"90919293", x"94979A9C", x"9D9F9F9E", x"9EA1A3A3", x"A3A1A1A3", x"A3A2A1A2",
									 -- x"A0A1A4A6", x"A6A3A3A4", x"A6A6A7A7", x"A7A8AAAC", x"A7ACAFB1", x"B2AFB0B6", x"B4B4B8BA", x"B7B8BAB8",
									 -- x"BBBCBCBC", x"BFC2C3C1", x"C2C4C5C4", x"C2C1C1C2", x"C8C7C7C9", x"CACBCAC9", x"C7C6C6C7", x"C6C5C5C7",
									 -- x"C4C2C1C2", x"C1C1C2C4", x"C1C1C0BF", x"BEBEBEBF", x"BFBCBBBB", x"B9B5B5B9", x"B7B4B6B8", x"B3AEABA7",
									 -- x"A4A4A29E", x"9D9E9D9A", x"98989794", x"918E8C8C", x"8A878585", x"827E7B7B", x"7B787778", x"78747171",
									 -- x"88878688", x"89888787", x"8A8A8A8A", x"8A8B8B8B", x"8C919396", x"9C9C9BA2", x"A2A2A1A2", x"A3A3A19F",
									 -- x"9D9B9999", x"9A989490", x"8F90908E", x"8B89898B", x"89888786", x"85848280", x"83848584", x"827F7E7D",
									 -- x"7C7C7A77", x"77777776", x"75797877", x"78767476", x"76767778", x"7B7E8081", x"83838586", x"88898888",
									 -- x"8C8A8889", x"88878788", x"8A898889", x"8A8A8A89", x"8B898888", x"88888989", x"8B8C8D8D", x"8E8E8E8F",
									 -- x"93919599", x"989A9FA1", x"A2A2A1A1", x"A09F9E9D", x"A1A09F9E", x"9E9D9C9B", x"9A9C9EA1", x"A3A5A7A9",
									 -- x"A9ABADAD", x"ADAEADAA", x"AEADACAD", x"AEAFAFAF", x"B3B1B0B1", x"B2B2B3B6", x"B5B4B5B8", x"BABABBBC",
									 -- x"BDBEBFC0", x"C1C2C3C3", x"C6C7C7C8", x"C9C9CACA", x"CCCBCBCD", x"CDCCCED1", x"CFD1D1CF", x"CECDCBC9",
									 -- x"C8C9C9C8", x"C8C7C7C7", x"C8C8C8C9", x"CACBCCCC", x"CDCDCDCC", x"CBCBCCCD", x"CDCCCCCE", x"CECCCBCB",
									 -- x"CBCCCDCD", x"CECDCBC9", x"C8C5C5C6", x"C4C5C6C2", x"C0C0C1C2", x"C4C5C5C5", x"C7CACDCF", x"D1D4D5D4",
									 -- x"D4D8DCDF", x"E0DFDFDF", x"E1E0DEDD", x"DDDFE1E2", x"E1E4E7E8", x"E8E7E7E7", x"E8EAEAE8", x"E6E6E7E8",
									 -- x"EBEDEEEC", x"E9E7E8EA", x"E9EBEEEF", x"F0EFEEED", x"EFEEEDEC", x"ECECEDEE", x"EFEDECEB", x"EAE9E9EB",
									 -- x"E9E8E8E7", x"E7E6E4E2", x"E2E2E2E2", x"E0DEDDDD", x"DDDDDCDB", x"D8D5D1CE", x"CCC8C2BE", x"BCBAB7B4",
									 -- x"B5B3B1AE", x"ACA9A7A6", x"A5A19C99", x"9895908D", x"8C888380", x"7F7E7A77", x"74726E6A", x"66656463",
									 -- x"5F5F5C59", x"54525152", x"4D4D4A47", x"474B4B47", x"46474747", x"46464648", x"46464544", x"43424141",
									 -- x"3B404243", x"4646494F", x"4C4D4E4F", x"50515253", x"5555585D", x"5D5B5E65", x"62636569", x"6E727476",
									 -- x"767A7D80", x"8484868C", x"92929395", x"97999B9C", x"A0A1A09E", x"9EA0A2A3", x"A6A5A4A5", x"A5A5A5A5",
									 -- x"A5A5A5A6", x"A3A0A0A2", x"A5A6A7A9", x"AAAAABAC", x"ADAFAFB1", x"B3B1B0B4", x"B4B5BABD", x"BBBABCBA",
									 -- x"BBBBBCBD", x"C0C3C2C0", x"BFC1C2C2", x"C3C3C5C6", x"C9CACACA", x"C8C6C6C6", x"C5C5C6C8", x"C7C4C4C5",
									 -- x"C1C1C2C1", x"BFBEC0C4", x"C1BFBCBC", x"BDBEBDBC", x"B9B9B9B7", x"B5B5B4B4", x"B1AEB1B3", x"AEAAA7A1",
									 -- x"A3A3A19E", x"9C9B9997", x"98969391", x"908E8A87", x"86858383", x"817D7A78", x"74777774", x"72716E6B",
									 -- x"8C8A898B", x"8B898786", x"8C8C8C8C", x"8C8B8B8B", x"90929396", x"9A9A9CA1", x"A1A1A2A3", x"A4A3A2A1",
									 -- x"A19F9E9D", x"9C999592", x"8C8E8E8D", x"8B8A8B8C", x"87888888", x"87878582", x"80838583", x"807E7D7D",
									 -- x"79797775", x"75777673", x"73767674", x"75747376", x"73747474", x"787C7F7F", x"83848587", x"898A8B8B",
									 -- x"8E8B8889", x"8A898888", x"8A898A8C", x"8C8B8A8A", x"88888888", x"8788898A", x"8E909192", x"93939494",
									 -- x"9694989C", x"9B9EA4A6", x"A6A6A6A6", x"A5A5A4A4", x"A7A6A5A4", x"A4A3A2A1", x"9EA0A2A5", x"A6A8AAAB",
									 -- x"A9ACAEAE", x"AFB0AFAD", x"B0AFAEAF", x"B1B2B2B1", x"B0B0B1B3", x"B4B2B2B3", x"B6B5B5B7", x"B9B9BABB",
									 -- x"BDBDBFC1", x"C2C2C2C2", x"C6C7C8C8", x"C8C9C9CA", x"CCCACBCD", x"CDCCCDD1", x"CFD1D2D0", x"CECDCBC9",
									 -- x"C5C6C6C6", x"C5C5C5C6", x"C7C7C8C9", x"C9CACBCB", x"CDCCCCCC", x"CCCCCDCD", x"D0CECCCD", x"CCCAC9CA",
									 -- x"CACACACB", x"CCCDCAC6", x"C6C5C6C6", x"C3C4C5C0", x"C3C3C4C5", x"C7C8C9C9", x"C7C9CCCD", x"CFD2D2D2",
									 -- x"D5D7DADC", x"DCDCDCDD", x"DEDDDCDC", x"DDDEE0E1", x"E0E2E5E6", x"E6E6E6E7", x"E7E8E9E7", x"E5E6E7E8",
									 -- x"EAECEDEB", x"E7E5E6E8", x"E7E8EBED", x"EEEFEFEE", x"EDECECEB", x"ECEDEEEF", x"EEEDEBEA", x"E9E9EAEB",
									 -- x"EAEAE9E8", x"E7E4E2E0", x"E3E2E3E3", x"E1DEDCDC", x"DCDAD8D6", x"D4D1CFCD", x"CAC6C0BE", x"BDBBB7B4",
									 -- x"B2AEAAA9", x"A8A7A5A4", x"9F9C9997", x"9694908D", x"8C89837E", x"7C7B7977", x"75736E69", x"66666461",
									 -- x"5F605F5B", x"55525153", x"504E4A47", x"47494845", x"47484848", x"47464647", x"43454646", x"45444444",
									 -- x"41444345", x"4848484D", x"4A4B4C4E", x"4F515355", x"5556585C", x"5D5C5F64", x"6565676C", x"6F727577",
									 -- x"7A7B7D82", x"898A888A", x"95949393", x"95989A9C", x"A2A2A1A0", x"9FA0A2A3", x"A5A4A3A3", x"A4A4A4A4",
									 -- x"A5A4A4A4", x"A2A0A1A4", x"A5A6A8A9", x"A9A9A9A9", x"AFB0AFB1", x"B6B5B3B6", x"B8B5B8BA", x"B8B9BBBB",
									 -- x"BABBBCBC", x"BFC1C0BE", x"C0C0C0C0", x"C1C2C4C5", x"C6C7C8C7", x"C5C3C3C3", x"C5C5C6C7", x"C6C2C1C1",
									 -- x"BFBFC0C0", x"BDBBBDC1", x"BFBCB9B9", x"BBBCBAB8", x"B5B6B7B6", x"B6B5B2AF", x"AEAAAAAB", x"A8A7A6A2",
									 -- x"A2A09E9D", x"9B979494", x"95928E8D", x"8D8C8783", x"8382807F", x"7E7B7876", x"73767570", x"6D6E6B67",
									 -- x"8F8D8D8F", x"918F8C8B", x"8E8D8C8B", x"8B8C8E8E", x"93919396", x"96989EA0", x"A1A2A3A4", x"A3A3A3A3",
									 -- x"A6A5A3A1", x"9E9B9794", x"8F8E8E8D", x"8D8C8B89", x"86888888", x"88898784", x"7F828482", x"807F7E7C",
									 -- x"75777877", x"76757472", x"73777674", x"75747377", x"73747475", x"787D7F7E", x"82838687", x"88898C8D",
									 -- x"8E8C8B8C", x"8B8A8889", x"8A898A8C", x"8D8B8A8B", x"86888A8A", x"89898B8E", x"90929596", x"97989A9B",
									 -- x"9B9A9EA3", x"A2A5AAAC", x"A9AAAAAB", x"ABABACAC", x"ADABAAA9", x"A9A9A9A8", x"A7A8AAAB", x"ACADAEAE",
									 -- x"AEB0B2B2", x"B3B4B3B1", x"B2B1B1B3", x"B5B7B6B5", x"B3B2B3B5", x"B5B3B2B3", x"B6B4B3B5", x"B8B9BABC",
									 -- x"BCBDBEC0", x"C1C1C2C2", x"C4C5C7C8", x"C8C8C9CA", x"CBC9CACD", x"CECCCED2", x"D0D2D3D1", x"CFCDCBC8",
									 -- x"C4C5C5C5", x"C4C4C5C6", x"C6C7C8C8", x"C9C9C9C9", x"CACACACB", x"CCCDCDCD", x"D0CDCBCB", x"CAC9C9C9",
									 -- x"CACCCCCB", x"CBCBC8C5", x"C5C5C7C6", x"C2C3C4C0", x"C0C1C2C2", x"C2C3C5C7", x"C7C9CBCB", x"CDD0D1D0",
									 -- x"D5D6D8D9", x"D9D9DADB", x"DADADBDB", x"DCDEDFDF", x"E1E2E3E3", x"E3E4E6E8", x"E7E8E7E5", x"E4E6E8E7",
									 -- x"EAEBECEA", x"E7E5E6E8", x"E7E7E9EA", x"ECEEEEEE", x"EBEBEBEC", x"ECEDEEEE", x"EBEBEAE9", x"E8E9E9E9",
									 -- x"E8E7E7E6", x"E4E2DFDD", x"DEDEE0E2", x"E0DCDADA", x"D8D7D5D3", x"D1CFCCCB", x"C6C3C0BE", x"BDBBB7B5",
									 -- x"AFABA7A6", x"A5A3A2A3", x"9C9A9895", x"93908D8B", x"8886827D", x"7A797876", x"76736E69", x"6868635E",
									 -- x"5F5F5E5A", x"56535252", x"514C4948", x"49484645", x"47474747", x"47464645", x"43444647", x"47464443",
									 -- x"47454244", x"4B4C494A", x"484A4D50", x"51525455", x"5456585A", x"5C5E6163", x"68686B6E", x"6F707478",
									 -- x"797C7E83", x"8A8B8A8E", x"94939294", x"979A9B9A", x"A1A1A1A1", x"A1A0A1A2", x"A0A0A0A1", x"A2A2A1A1",
									 -- x"A2A1A2A2", x"A2A1A3A6", x"A5A6A8A8", x"A7A7A8A9", x"ABADADB2", x"B8B7B5B7", x"B9B4B5B7", x"B6B7BABA",
									 -- x"BBBCBCBB", x"BCBEBFBD", x"C2C0BEBE", x"BEC0C1C1", x"C2C3C3C3", x"C3C2C2C2", x"C3C2C3C4", x"C3C0BFBF",
									 -- x"BFBDBCBC", x"BCBABABB", x"BBB9B7B8", x"B9B9B8B6", x"B6B2B1B4", x"B5B2AEAD", x"AEA9A7A5", x"A2A3A4A0",
									 -- x"9F9A999A", x"97919093", x"8F8D8B8A", x"89878481", x"817E7B79", x"79787573", x"7272716F", x"6E6C6965",
									 -- x"95939295", x"9593908E", x"8D8C8A8A", x"8B8D9092", x"928E9195", x"92979FA1", x"A5A6A7A7", x"A6A5A5A6",
									 -- x"A6A6A5A4", x"A19E9B99", x"97939090", x"92908C88", x"86888887", x"87888784", x"83858582", x"807F7C78",
									 -- x"73777B7A", x"77757372", x"74777674", x"7575757A", x"76777777", x"7B7F807E", x"80828586", x"86888B8E",
									 -- x"8D8D8E8E", x"8D8A898A", x"8988898C", x"8D8B8B8C", x"86898D8D", x"8C8C8F92", x"8F929698", x"9A9B9D9F",
									 -- x"A1A0A5AA", x"A9ABAFB0", x"B2B2B2B1", x"B0AFB0B0", x"B1AFADAC", x"ACADAEAE", x"AEAFB1B1", x"B1B1B1B1",
									 -- x"B4B6B7B6", x"B6B7B6B4", x"B3B2B3B5", x"B9BBBAB9", x"BBB9B7B7", x"B6B5B5B7", x"B5B2B1B4", x"B7B9BBBD",
									 -- x"BCBDBDBE", x"BFC0C1C2", x"C2C4C6C7", x"C7C8C9CA", x"CBC8C9CD", x"CECCCED3", x"D0D2D3D1", x"CFCDC9C6",
									 -- x"C6C6C6C6", x"C4C4C6C7", x"C6C6C7C8", x"C9C9C8C8", x"C8C8C9CA", x"CBCCCDCD", x"CFCBC9C9", x"C9C9C9CB",
									 -- x"CACDCECC", x"C9C9C7C5", x"C4C5C8C6", x"C1C2C3BF", x"C0C2C2C1", x"C0C1C4C7", x"C7C8CACA", x"CCCFD1D0",
									 -- x"D2D3D4D4", x"D4D5D7D9", x"D7D8DADB", x"DDDDDDDD", x"E1E1E1E0", x"E0E3E7EA", x"E8E9E7E4", x"E4E7E8E7",
									 -- x"EBEBEBEA", x"E7E6E7E8", x"E8E8E8E9", x"EAECECED", x"EBEBECEC", x"EDECECEB", x"E9EAEAE9", x"E8E8E7E6",
									 -- x"E4E4E3E3", x"E2E0DDDB", x"D9DADCDF", x"DEDAD7D7", x"D3D2D0CE", x"CDCBC9C7", x"C4C3C1BD", x"B9B4B1AF",
									 -- x"ADA8A5A3", x"A19E9E9F", x"9C9B9894", x"908C8987", x"8283817C", x"79787776", x"73716C68", x"6867615A",
									 -- x"5C5B5957", x"5552504E", x"4F4A474A", x"4B494747", x"46464646", x"47474544", x"44444547", x"48474441",
									 -- x"42454648", x"4A484A51", x"4D4F5254", x"53525151", x"5457595B", x"5F636665", x"68686A6D", x"6D6D7075",
									 -- x"737A7F82", x"85848992", x"90919398", x"9C9D9C9A", x"9C9D9E9F", x"9F9E9E9F", x"9FA0A1A2", x"A3A3A2A0",
									 -- x"A4A3A3A4", x"A3A1A3A5", x"A5A7A8A7", x"A6A6A9AB", x"A9ACAEB2", x"B7B5B2B4", x"B9B4B5B9", x"B9BABCBA",
									 -- x"BCBDBCBA", x"BABCBEBD", x"BFBDBBBB", x"BDC0C2C2", x"C4C3C1C1", x"C2C2C1BF", x"C0BFC0C1", x"C0BEBEC0",
									 -- x"BFBAB8B9", x"BBB9B7B5", x"B8B8B8B8", x"B8B7B7B6", x"B9AEAAAE", x"B0ABA9AD", x"ABA6A4A2", x"9E9F9E9A",
									 -- x"9C959396", x"948D8D93", x"89898887", x"86848180", x"7F7C7875", x"74747271", x"6E6A6A70", x"716C6562",
									 -- x"95969695", x"92919192", x"8C8A8B8E", x"8F8E8F90", x"92919293", x"9395999E", x"A6A6A6A7", x"A6A5A6A7",
									 -- x"A6A9A9A6", x"A5A39E96", x"93949491", x"8F8E8C89", x"89888584", x"86898986", x"88878583", x"817E7B7A",
									 -- x"7A797776", x"75757576", x"78787674", x"75787775", x"7573777C", x"7B7B7F7F", x"80808386", x"87858789",
									 -- x"8E909495", x"918C8C8F", x"888A8D8E", x"8E8C8A89", x"8C8C8D8F", x"8F8F9195", x"92969999", x"9DA2A3A0",
									 -- x"A6A8ABAC", x"AEB1B6BA", x"B6B7B7B5", x"B3B3B4B5", x"B2B2B2B1", x"B1B1B3B4", x"B2B2B3B5", x"B8BABBBB",
									 -- x"B8BCBEBE", x"BEBFBFBE", x"BABBBBBB", x"BBBBBBBB", x"BCBDBCBB", x"B8B7B6B7", x"B6B4B4B5", x"B7BABCBC",
									 -- x"BBBDBEBE", x"BFC2C3C4", x"C2C5C7C8", x"C7C7C8C9", x"C7C7C9CC", x"CDCDCFD2", x"D3D3D2D1", x"CFCCC8C6",
									 -- x"C5C5C6C7", x"C6C4C5C7", x"C5C7C7C5", x"C5C6C5C4", x"C5C6C7C9", x"CACBCBCB", x"CCCBCAC9", x"CACBCCCC",
									 -- x"CDCBC9C8", x"C8C8C6C5", x"C6C5C3C2", x"C2C4C5C6", x"C4C2C1C2", x"C3C2C1C2", x"C8C9CBCC", x"CDCECFD0",
									 -- x"CDD0D4D6", x"D6D7D6D5", x"D4D7D9D9", x"DADCDDDD", x"DDDFE2E4", x"E4E4E5E6", x"E7E7E6E5", x"E5E6E7E8",
									 -- x"E8E8E9E8", x"E7E7E7E7", x"E6E8E9EA", x"EAEAEAEA", x"E8EAEAE9", x"E9EBEAE7", x"E7E7E7E7", x"E7E7E5E4",
									 -- x"E2E4E4E2", x"DFDDDEDF", x"DCDCDCDA", x"D8D7D6D5", x"D2D0CECD", x"CDCBC8C6", x"C5C0BCBB", x"B9B5B0AE",
									 -- x"AAA8A5A2", x"9F9D9A99", x"96979592", x"8E8C8A88", x"83827F7B", x"78777676", x"77706A68", x"6764605F",
									 -- x"59595855", x"54555552", x"4F4E4B47", x"45464A4D", x"48474646", x"46454342", x"46454445", x"46454341",
									 -- x"42434446", x"4545494D", x"4B4E5150", x"4F4E4F50", x"51595B5B", x"5E616366", x"6F6C696B", x"6D6F7275",
									 -- x"77797D80", x"8284898F", x"8B91989B", x"9B9DA1A4", x"9C9EA29E", x"A49D9E9E", x"A19E9C9F", x"A1A1A2A3",
									 -- x"A3A5A5A3", x"A3A5A3A1", x"A5A3A3A4", x"A5A5A7A9", x"A7AAACAC", x"AFB3B5B3", x"B7B5B6B8", x"BAB9B9BB",
									 -- x"BDBDBCBC", x"BCBCBCBC", x"B9BCBFC1", x"C0BEBEBE", x"C0BFBEBE", x"BFBEBEBE", x"BBC0BDBA", x"BCB9B8BF",
									 -- x"BAB9BABB", x"B8B4B5B8", x"B5B7B4AE", x"AFB3B0A9", x"ACAFB1B0", x"ACA8A6A6", x"A0A3A4A0", x"9B9E9D95",
									 -- x"98979692", x"8E8B8A8A", x"89868585", x"837E7A79", x"7C777372", x"72707070", x"6E6E6B66", x"66696965",
									 -- x"96969595", x"94949495", x"93908F91", x"93919090", x"91909192", x"9394979A", x"A2A3A5A6", x"A6A7A7A7",
									 -- x"A7A9A9A6", x"A4A39E97", x"97979490", x"8D8C8A87", x"89888786", x"888A8986", x"85848281", x"807E7C7A",
									 -- x"79797877", x"76757575", x"75757573", x"74777775", x"77777C80", x"7D7D8183", x"82828588", x"89888A8D",
									 -- x"90909396", x"96939192", x"8D8C8C8B", x"8A8B8C8D", x"8E8E8F90", x"90919498", x"999B9D9F", x"A1A4A5A4",
									 -- x"A9ABAEB0", x"B3B6BBBE", x"BCBCBAB9", x"B7B6B7B7", x"B9B9B8B7", x"B5B5B5B6", x"B5B6B7B9", x"BCBEBFC0",
									 -- x"BDC0C1C0", x"C0C1C1C1", x"BEBEBEBE", x"BEBEBEBD", x"BDBEBDBC", x"BAB9B9B9", x"B9B8B7B8", x"B9BBBBBB",
									 -- x"BCBEC0BF", x"C0C2C3C2", x"C3C5C7C8", x"C8C8C9CA", x"CACACBCD", x"CECDCED1", x"D2D2D2D2", x"D0CECBC9",
									 -- x"C6C5C6C7", x"C6C4C5C7", x"C5C7C7C6", x"C6C7C6C5", x"C5C5C6C7", x"C8C9CACB", x"CCCBCACA", x"CACACACA",
									 -- x"CBCAC9C8", x"C7C7C6C6", x"C4C4C3C3", x"C4C4C4C3", x"C3C1C1C2", x"C2C1C2C4", x"C8C9CBCC", x"CECFCFD0",
									 -- x"CECFD2D3", x"D4D5D6D7", x"D7D9DAD9", x"DADBDCDC", x"DEDFE1E2", x"E2E3E4E6", x"E5E5E4E4", x"E4E5E5E6",
									 -- x"E5E5E6E6", x"E5E6E7E8", x"E6E7E8E9", x"E9E8E9E9", x"E9EAEAE9", x"E9EAE9E6", x"E6E6E6E6", x"E6E5E4E3",
									 -- x"E0E2E2E0", x"DDDBDBDD", x"DDDCDBD9", x"D7D5D5D5", x"D2D0CECC", x"CBC9C6C4", x"C0BEBCBB", x"B7B2AEAD",
									 -- x"A9A8A5A2", x"A09E9D9C", x"97989793", x"908E8B89", x"8784807E", x"7C797674", x"6F6F706E", x"69626061",
									 -- x"5E5E5C59", x"58585653", x"4F4F4E4C", x"4A494A4C", x"47474645", x"43434343", x"48464444", x"44454544",
									 -- x"45454648", x"48484A4D", x"4E4F5051", x"51525353", x"545B5C5B", x"5E606165", x"68696C6F", x"71717377",
									 -- x"7C7D8083", x"8384888C", x"8E929698", x"9A9C9FA2", x"9C9E9B9C", x"9EA09FA1", x"A29F9EA0", x"A1A0A1A3",
									 -- x"A1A2A2A0", x"9FA09F9D", x"A5A4A4A5", x"A4A4A6A9", x"AAACADAE", x"B0B4B5B4", x"B9B6B6B9", x"BBBBBBBB",
									 -- x"BBBBBBBC", x"BCBCBDBE", x"BCBDBEBE", x"BEBDBDBD", x"BEBDBCBB", x"BABABABA", x"B9BDBDBB", x"B9B7B7BB",
									 -- x"B6B6B6B7", x"B5B4B4B6", x"B3B2B0AF", x"AFAFACA9", x"A9ABADAC", x"A8A5A4A5", x"A3A09E9C", x"9897958F",
									 -- x"9494928F", x"8B888787", x"85838181", x"7F7A7777", x"79747070", x"706E6E6E", x"6B6B6863", x"63656562",
									 -- x"9B999796", x"96959594", x"93919092", x"95949393", x"92909193", x"95959597", x"9B9FA2A3", x"A4A8A9A8",
									 -- x"A9ABAAA8", x"A7A7A39E", x"9E9B9691", x"8F8E8C89", x"89898887", x"898A8784", x"82817F7E", x"7E7D7C7B",
									 -- x"79797979", x"78777675", x"74757574", x"74757676", x"78797F82", x"7D7D8183", x"8385878A", x"8B8B8E91",
									 -- x"91909296", x"99989593", x"92908E8C", x"8C8D8F91", x"90909192", x"9393979A", x"9F9E9FA2", x"A4A4A6A7",
									 -- x"ACAEB2B5", x"B8BCC0C3", x"C2C0BEBC", x"BBBBBBBB", x"BEBEBEBC", x"BBB9B8B8", x"B9B9BABC", x"C0C2C4C4",
									 -- x"C2C4C4C3", x"C2C3C4C3", x"C3C2C1C2", x"C3C3C2C1", x"C0BFBFBD", x"BCBBBCBC", x"B9B8B8B9", x"BABABABA",
									 -- x"BBBEC0C1", x"C1C3C3C2", x"C3C5C7C9", x"C9C9CBCC", x"CCCCCCCE", x"CECDCFD1", x"D2D2D3D2", x"D1CFCCCA",
									 -- x"C7C6C6C7", x"C6C5C5C7", x"C5C6C7C6", x"C6C7C7C6", x"C6C6C6C6", x"C7C8CACB", x"CCCBCBCB", x"CBCBCAC9",
									 -- x"C8C9C9C8", x"C6C5C6C7", x"C1C2C3C4", x"C5C4C2C1", x"C2C1C1C2", x"C1C0C2C6", x"C8C9CBCD", x"CFD0CFCF",
									 -- x"CFD0D1D2", x"D3D4D5D7", x"D8D9DAD8", x"D8DADBDA", x"DDDEDFDF", x"DFE0E2E5", x"E2E2E2E2", x"E2E2E3E3",
									 -- x"E2E2E2E2", x"E3E4E6E7", x"E5E6E7E7", x"E7E6E7E7", x"E8E8E8E7", x"E7E8E6E4", x"E5E5E4E4", x"E4E3E2E0",
									 -- x"DEDFDFDD", x"DBD9D8D9", x"DAD9D7D6", x"D4D4D3D4", x"D1CFCCCA", x"C9C7C4C2", x"BDBCBCBB", x"B6B0ADAC",
									 -- x"A9A7A5A2", x"9F9D9C9C", x"9292918E", x"8B898683", x"84807C7B", x"7A78736F", x"6D6F716F", x"6A636162",
									 -- x"5F5F5D5A", x"58585653", x"4F4F4E4C", x"4A4A4A4B", x"47474744", x"41414345", x"44454647", x"47474645",
									 -- x"4646474A", x"4B4A4A4C", x"4D4C4C4D", x"4F505050", x"54595A5A", x"5E616468", x"65696E72", x"7271757A",
									 -- x"797B7F83", x"85878B90", x"94949597", x"9A9D9FA0", x"9D9F979B", x"999F999D", x"9E9D9D9E", x"9D9D9EA0",
									 -- x"A1A3A3A1", x"A0A0A1A1", x"A4A4A5A5", x"A4A3A6A9", x"ACAEAEAF", x"B0B3B5B5", x"B7B5B5B8", x"BBBCBBBB",
									 -- x"B9BABBBB", x"BABABBBC", x"BDBCBBBA", x"BBBCBCBC", x"BABDBCB8", x"B6B8B9B9", x"B6B8BBBB", x"B7B5B7B7",
									 -- x"B8B8B6B3", x"B2B2B2B0", x"AFADADAF", x"AEA9A7A8", x"A7A7A8A6", x"A3A1A0A0", x"9F979598", x"96949390",
									 -- x"8F8E8C8A", x"87848483", x"827F7D7C", x"7A787675", x"75716E6D", x"6C6B6A6A", x"65666360", x"5F61615F",
									 -- x"9D9A9797", x"98989693", x"93939495", x"96969696", x"95929295", x"97989797", x"979C9F9F", x"A1A7AAA9",
									 -- x"ABACABAA", x"AAABA9A5", x"A29E9792", x"9192908D", x"88888785", x"86868481", x"807E7D7C", x"7C7B7A7A",
									 -- x"7A7A7A7A", x"79787777", x"76777876", x"75757676", x"79797F81", x"7E7E8182", x"8586898B", x"8C8E9194",
									 -- x"91909195", x"99999693", x"92919090", x"90909090", x"91929495", x"9697999B", x"A19FA1A5", x"A7A6A8AC",
									 -- x"AFB2B6BA", x"BDC0C3C5", x"C5C3BFBE", x"BEBFBFBF", x"BEBFBFBF", x"BEBCBBBB", x"BABABBBD", x"C0C3C5C6",
									 -- x"C4C6C7C6", x"C5C6C6C4", x"C6C5C5C6", x"C8C8C7C6", x"C3C2C1C0", x"BEBDBDBE", x"BABABABA", x"BABBBCBC",
									 -- x"BBBEC1C1", x"C2C3C3C2", x"C3C5C7C9", x"CACCCDCE", x"CBCBCBCC", x"CDCECFD1", x"D2D3D3D2", x"D0CDCBCA",
									 -- x"C8C7C7C7", x"C7C5C5C7", x"C5C7C7C6", x"C6C7C6C5", x"C6C6C6C7", x"C7C8C9CA", x"CAC9C9C9", x"C9C9C7C6",
									 -- x"C8C7C6C6", x"C5C4C4C4", x"C0C0C1C3", x"C4C3C2C1", x"C4C3C3C3", x"C1C0C2C6", x"C9CACBCE", x"D0D0CFCE",
									 -- x"D1D1D1D2", x"D3D3D4D6", x"D6D8D7D6", x"D6D8D9D9", x"DBDCDDDD", x"DCDDE0E2", x"E0E0E0E0", x"E0E0E0E0",
									 -- x"E1E1E1E0", x"E0E1E3E5", x"E3E4E4E5", x"E4E4E5E5", x"E5E6E5E5", x"E6E5E4E3", x"E5E4E4E3", x"E3E2E0DF",
									 -- x"DDDDDCDB", x"D9D7D6D5", x"D4D3D3D2", x"D2D2D2D1", x"CFCDCAC8", x"C7C5C3C1", x"BBBAB9B7", x"B3AFACAA",
									 -- x"A9A8A5A1", x"9D9A9998", x"9393908C", x"8A898885", x"807E7B79", x"79787471", x"73706D6B", x"6A676563",
									 -- x"5E5E5C5A", x"59575554", x"514F4B48", x"47484A4B", x"48484644", x"43434445", x"44454546", x"4748494A",
									 -- x"4645474A", x"4C4B4A4A", x"51505051", x"52525253", x"55595A5A", x"5F62656A", x"6A6C6F70", x"7071767C",
									 -- x"76787C82", x"85888D92", x"95939295", x"999D9D9C", x"9DA09B9D", x"9C9E9A9C", x"9B9C9D9C", x"9B9B9D9F",
									 -- x"A2A4A5A4", x"A2A2A4A6", x"A2A3A5A7", x"A5A4A6AA", x"ACADAEAE", x"AFB2B4B5", x"B2B2B3B5", x"B8B9BABB",
									 -- x"B9BABBBA", x"B8B7B8B9", x"BBB9B7B7", x"B9BABBBA", x"B6BABAB5", x"B3B6B9B8", x"B5B2B7BA", x"B6B6B8B3",
									 -- x"B6B7B4AE", x"ADAFAEAB", x"ABABACAE", x"ABA6A4A5", x"A5A5A4A2", x"9F9D9B9A", x"98939295", x"94949390",
									 -- x"8A898785", x"83818080", x"7D7B7876", x"75747372", x"716F6C6A", x"69676666", x"6162605D", x"5D5E5F5D",
									 -- x"9A989698", x"9B9C9A98", x"999B9C9A", x"98979798", x"98959396", x"999A9A9A", x"969A9B9B", x"9EA4A8A8",
									 -- x"ABABAAAA", x"AAABA9A6", x"A39F9892", x"9192908D", x"87868481", x"8182807E", x"7F7E7C7B", x"7B7A7978",
									 -- x"7B7A7A79", x"78787878", x"77787877", x"76757678", x"7B7A7E81", x"80828481", x"85888A8B", x"8D8F9294",
									 -- x"92939496", x"97979593", x"90908F90", x"9090908F", x"91949798", x"999A9B9C", x"A5A4A6AA", x"ABAAADB1",
									 -- x"B5B8BCC0", x"C3C5C6C6", x"C7C4C1C0", x"C0C1C1C0", x"C0C1C1C1", x"C0BEBDBD", x"BCBCBCBE", x"C1C4C5C6",
									 -- x"C6C8CACA", x"CACAC9C6", x"C8C7C7C8", x"CACCCCCC", x"C8C7C5C3", x"C1C0BFBE", x"BFBFBEBE", x"BEBEBFC0",
									 -- x"BDC0C2C2", x"C2C3C3C2", x"C4C5C7C9", x"CBCDCFD0", x"CCCBCBCB", x"CCCDCECE", x"D0D1D2D1", x"CFCCCBCB",
									 -- x"CAC8C7C8", x"C8C6C6C7", x"C6C7C7C6", x"C5C6C5C4", x"C5C5C6C7", x"C7C7C7C7", x"C6C6C6C6", x"C7C6C4C3",
									 -- x"C8C6C3C3", x"C4C4C2BF", x"C0BFBFBF", x"C1C2C3C3", x"C3C3C3C3", x"C1C1C4C8", x"CACBCDCE", x"D0D0CFCD",
									 -- x"D1D1D2D4", x"D5D4D5D7", x"D7D8D7D5", x"D5D7D8D8", x"DADCDDDD", x"DDDDDEE0", x"DEDEDEDE", x"DEDEDFDF",
									 -- x"DFDFDFDF", x"DEDFE1E3", x"E1E2E2E2", x"E2E2E3E4", x"E4E4E4E5", x"E5E5E4E4", x"E5E4E3E3", x"E2E1DFDE",
									 -- x"DCDBDAD9", x"D8D6D4D2", x"D1D0D0D1", x"D1D1CFCD", x"CDCBC9C7", x"C5C3C0BE", x"BAB8B5B2", x"B0AEABA8",
									 -- x"A9A8A5A1", x"9C989797", x"9594908B", x"898A8987", x"82817F7D", x"7C7A7978", x"74716D6A", x"69686764",
									 -- x"615F5E5D", x"5B595655", x"52504C49", x"48494A4B", x"4A484646", x"48484644", x"4A474442", x"43474C4F",
									 -- x"4948494B", x"4C4A4948", x"50505355", x"54525356", x"5B5D5C5C", x"5F606267", x"6E6D6D6F", x"7073777C",
									 -- x"7A7B7F83", x"86878B8E", x"918F8F92", x"979A9A98", x"9B9EA09C", x"A19EA1A4", x"9FA0A09F", x"9E9D9E9F",
									 -- x"A0A1A2A2", x"A0A0A2A5", x"A0A2A5A7", x"A7A6A7AA", x"ACACADAE", x"AFB1B3B6", x"B1B3B6B6", x"B6B7B9BA",
									 -- x"BABBBBBA", x"B8B7B6B7", x"BAB8B7B7", x"B8B9B8B7", x"B2B5B5B1", x"AFB1B4B4", x"B3AEB1B5", x"B3B4B3AC",
									 -- x"ADAEACA8", x"A8ABABA9", x"A7ABADAA", x"A6A4A2A0", x"A2A1A09F", x"9D9A9896", x"94939493", x"8F8F8E89",
									 -- x"86858381", x"807E7D7C", x"77767371", x"70706F6E", x"6D6C6A68", x"67666563", x"61615F5D", x"5B5B5B5B",
									 -- x"9E9C9A9B", x"9D9D9B99", x"9A9C9D9C", x"99999A9A", x"99969598", x"9A9B9A9A", x"9899999A", x"9C9FA3A6",
									 -- x"ADACABAA", x"ABAAA8A6", x"A5A29C96", x"94928F8C", x"8786837F", x"7E7E7E7C", x"7F7E7C7B", x"7A7A7A79",
									 -- x"7B7A7978", x"78777778", x"78777677", x"7776787A", x"7A7A7E81", x"82858681", x"878A8C8D", x"8E919394",
									 -- x"95979897", x"97989795", x"93918F8F", x"91929393", x"93979A9B", x"9C9E9F9F", x"A8A8ABAD", x"AEAEB0B3",
									 -- x"BCBEC2C6", x"C9CAC9C8", x"C9C8C5C3", x"C3C3C3C3", x"C5C5C5C4", x"C2C0BFBE", x"BEBEBEC0", x"C3C5C7C8",
									 -- x"CACCCECF", x"CFCFCCC9", x"CACACACA", x"CCCED0D1", x"CECDCAC8", x"C7C4C2C0", x"C2C2C2C1", x"C0BFC0C0",
									 -- x"C0C3C4C3", x"C3C4C4C3", x"C6C6C8C9", x"CBCDCFD0", x"CECECCCB", x"CBCDCDCC", x"CECFD1D0", x"CFCDCDCE",
									 -- x"CCCAC8C9", x"C9C8C7C8", x"C7C8C8C6", x"C6C6C5C4", x"C3C4C4C5", x"C5C5C4C4", x"C5C6C6C7", x"C7C7C6C5",
									 -- x"C8C5C1C1", x"C3C3C0BD", x"BFBEBEBE", x"BFC1C2C2", x"C1C0C1C2", x"C3C3C6C9", x"CACCCECF", x"CFCFCFCF",
									 -- x"D0CFD2D5", x"D7D5D6DA", x"D9DAD9D6", x"D5D6D8D7", x"DADCDDDE", x"DDDDDDDE", x"DDDCDCDC", x"DCDDDDDD",
									 -- x"DDDDDEDD", x"DDDEE0E1", x"DFE0E0E0", x"E0E1E2E3", x"E4E3E4E5", x"E6E5E5E5", x"E4E3E3E2", x"E2E1DFDE",
									 -- x"DBDAD9D8", x"D7D5D2D0", x"D1D1D0D0", x"D0CFCBC9", x"CBC9C7C5", x"C3C0BDBA", x"BCB9B5B2", x"B1B1ADAA",
									 -- x"A7A7A5A2", x"9D999898", x"95938E89", x"88898987", x"8483817E", x"7B797877", x"7072716D", x"69676564",
									 -- x"62605E5D", x"5B585554", x"53514F4E", x"4D4C4B4A", x"4A484749", x"4B4C4946", x"48474646", x"48494949",
									 -- x"4C4B4C4D", x"4C4A494A", x"4C4D5155", x"54525458", x"5C5D5C5D", x"60616368", x"6C6A6B6F", x"73757779",
									 -- x"7C7D8084", x"87888B8D", x"8E8E9093", x"989A9A99", x"9B9DA098", x"9E99A0A5", x"A1A2A2A0", x"9E9E9E9D",
									 -- x"9E9E9F9F", x"9E9D9EA1", x"A0A0A2A5", x"A7A6A7A9", x"ACACAEAF", x"B0B0B3B6", x"B4B6B8B6", x"B5B5B6B7",
									 -- x"B8B8B8B8", x"B8B7B7B6", x"B8B8B8B7", x"B7B6B5B4", x"B3B3B2B0", x"AEADAEB0", x"B0ACABAE", x"AFAFACA6",
									 -- x"ABABA9A6", x"A5A6A7A7", x"A5A9A9A5", x"A2A19F9C", x"9D9B9A99", x"99989593", x"8E8F908E", x"88898882",
									 -- x"82817F7D", x"7C7B7978", x"74747270", x"6F6F6D6B", x"67676765", x"64646362", x"61605F5C", x"59575757",
									 -- x"A7A4A09E", x"9D9D9B9A", x"9B9C9C9B", x"9C9E9D9B", x"9A98989B", x"9C9B9A9A", x"9B98989A", x"9B9A9DA2",
									 -- x"ABAAA9AA", x"ABAAA8A6", x"A7A5A19B", x"96938F8B", x"89888580", x"7E7E7E7C", x"7E7D7B7B", x"7B7C7C7C",
									 -- x"7B7B7B7B", x"7B7A7979", x"7B787677", x"7878797C", x"797B8083", x"83878985", x"898D8F8F", x"90929494",
									 -- x"98999998", x"989A9997", x"96949292", x"94969797", x"989C9E9E", x"9FA2A4A4", x"A9ADB0B1", x"B2B4B7B8",
									 -- x"C0C3C7CB", x"CDCDCCCA", x"CACAC9C8", x"C8C8C9CA", x"C9C9C9C7", x"C5C2C1C0", x"C0C0C0C2", x"C5C8CACB",
									 -- x"CFD0D1D1", x"D2D2CFCB", x"CCCCCCCC", x"CCCED2D5", x"D4D2D0CF", x"CDCAC7C4", x"C2C3C5C5", x"C3C2C1C1",
									 -- x"C3C4C5C3", x"C4C6C7C7", x"C8C8C9CA", x"CBCCCDCD", x"D1D0CECC", x"CCCECECD", x"CFD0D2D2", x"D0CFCFD0",
									 -- x"CECBC9CA", x"CAC9C8C9", x"C8C9C9C7", x"C7C8C7C5", x"C3C3C3C3", x"C3C3C3C3", x"C6C6C6C7", x"C8C9C8C7",
									 -- x"C7C4C1C1", x"C3C3C1BE", x"BEBEBEBF", x"C0C0C0BF", x"BFBEBFC1", x"C3C4C6C8", x"C9CCCFCF", x"CECED0D2",
									 -- x"D2D0D2D6", x"D7D5D6DA", x"D9DAD9D7", x"D5D7D7D7", x"D8DADBDB", x"DBDADBDC", x"DBDBDADA", x"DADBDCDC",
									 -- x"DCDDDDDD", x"DCDCDDDE", x"DEDEDFDF", x"DFE0E2E3", x"E4E2E3E5", x"E6E4E3E4", x"E3E2E2E1", x"E1E0DFDD",
									 -- x"DBD9D7D7", x"D7D5D1CE", x"D1CFCECD", x"CDCCC8C6", x"C6C5C4C3", x"C2BFBBB9", x"BABAB7B3", x"B1B1AEAB",
									 -- x"A5A5A5A2", x"9D9A9898", x"9795918D", x"8C8D8B89", x"83817F7D", x"7B787573", x"7172716D", x"6A686561",
									 -- x"605D5C5C", x"5A565352", x"52514F4D", x"4D4C4A49", x"4A49484A", x"4C4D4B49", x"45454649", x"4C4C4945",
									 -- x"4B4B4C4D", x"4C4B4C4F", x"52525459", x"5A595A5E", x"5A5B5B5D", x"6263656A", x"6B696B6F", x"73757778",
									 -- x"7C7C8084", x"87898B8D", x"8F919396", x"999B9C9D", x"9B9D9B98", x"99989A9F", x"9E9F9E9C", x"9C9D9C99",
									 -- x"9C9B9B9E", x"9F9E9EA0", x"A19F9FA1", x"A4A5A6A8", x"ABACAEB0", x"AFAEB0B4", x"B3B4B3B2", x"B2B4B3B1",
									 -- x"B4B3B3B4", x"B5B5B4B2", x"B3B4B5B5", x"B4B3B2B2", x"B4B1AFB0", x"AEABABAD", x"AAAAA8A8", x"ABAAA7A6",
									 -- x"ADABAAA8", x"A5A3A3A5", x"A4A3A2A1", x"9F9C9B9B", x"98969393", x"9393918F", x"8B878788", x"8583827E",
									 -- x"7F7D7B79", x"78777674", x"7171706E", x"6D6D6A67", x"63646462", x"60605F5E", x"5D5D5C59", x"56535353",
									 -- x"AAA7A29F", x"9E9E9F9F", x"A2A19E9D", x"9FA19E99", x"9B9A9C9E", x"9E9C9A9A", x"9C98989B", x"9B98999F",
									 -- x"A6A5A5A7", x"A8A8A7A6", x"A4A4A19B", x"96928E8A", x"8A898782", x"807F7E7D", x"7D7C7B7B", x"7C7D7E7E",
									 -- x"7D7E7E7F", x"7E7D7C7B", x"7F7B7879", x"7A797A7C", x"7B7E8587", x"868A8D8B", x"8B8F9291", x"92949594",
									 -- x"99999897", x"999C9B98", x"95939293", x"96979796", x"9C9FA1A0", x"A1A5A8A9", x"ABB1B5B6", x"B7BCBEBE",
									 -- x"C1C4C8CD", x"CFCFCCCA", x"CACBCCCC", x"CCCDCFD1", x"CBCBCAC8", x"C6C4C3C2", x"C0C0C0C2", x"C6C9CCCD",
									 -- x"D2D3D2D1", x"D2D2D0CC", x"CDCECECD", x"CCCED2D7", x"D7D6D4D3", x"D1CECAC8", x"C2C4C8C9", x"C8C6C4C4",
									 -- x"C3C4C5C4", x"C5C8CBCC", x"CBCACACA", x"CBCBCCCC", x"D1D1CFCD", x"CED1D1CF", x"D1D3D4D3", x"D1D0D0D1",
									 -- x"CFCCCACA", x"CAC9C9C9", x"C8C9CAC8", x"C8C9C8C7", x"C5C4C3C3", x"C2C3C3C4", x"C3C3C3C5", x"C6C7C7C7",
									 -- x"C5C4C3C2", x"C2C2C1C0", x"BDBDBFC1", x"C1C0BDBB", x"BFBDBEC1", x"C3C4C5C6", x"C8CBCFCF", x"CECED1D4",
									 -- x"D5D2D2D5", x"D5D3D4D8", x"D6D8D8D6", x"D5D7D8D7", x"D6D8D8D8", x"D7D7D8DA", x"DBDAD9D8", x"D9D9DBDB",
									 -- x"DDDDDDDC", x"DBDADADA", x"DDDEDEDE", x"DFE0E2E3", x"E3E1E1E3", x"E4E2E1E1", x"E2E1E1E1", x"E0E0DEDD",
									 -- x"DAD8D6D6", x"D6D4D0CD", x"CECCCACA", x"CAC9C7C4", x"C1C0C0C1", x"C1BFBCB9", x"B5B7B6B2", x"AEADABA8",
									 -- x"A3A4A4A1", x"9C989696", x"92908D8A", x"89898784", x"86838180", x"807D7874", x"77736D69", x"6B6C655E",
									 -- x"5E5C5B5B", x"5A565454", x"524F4B48", x"48484848", x"49494A4B", x"4C4C4C4B", x"4A454142", x"474C4D4C",
									 -- x"48494A4C", x"4C4C4F54", x"54515156", x"5958595C", x"5C5D5C5E", x"62626368", x"6C6A6B6E", x"71737679",
									 -- x"7D7D8084", x"8687888A", x"8F919496", x"98999C9E", x"979C989C", x"9A9E999E", x"9A9B9B9A", x"9B9D9C99",
									 -- x"9896989C", x"9F9F9FA1", x"A39F9C9E", x"A1A3A5A7", x"AAABADAF", x"AEACAEB1", x"AFAEACAC", x"AFB2B0AB",
									 -- x"B0AFAEAF", x"B2B2AFAC", x"ACAEB0B1", x"B0B0B0B1", x"B1ABAAAD", x"ADA8A7AB", x"A5A9A7A6", x"AAA9A6AA",
									 -- x"A8A7A6A7", x"A4A1A2A7", x"A49E9C9F", x"9E98979B", x"97938F8E", x"8E8E8D8B", x"8E848185", x"837E7C7B",
									 -- x"7C7A7877", x"76757371", x"6B6D6C6A", x"69686561", x"62646360", x"5D5D5B59", x"59595856", x"54515152",
									 -- x"ADABA7A4", x"A19F9F9F", x"9F9F9E9E", x"9F9F9F9E", x"A09E9C9C", x"9D9E9D9C", x"9B9A9A9A", x"9B9C9D9D",
									 -- x"A3A4A7A9", x"AAAAA8A7", x"A29F9C9A", x"9995908C", x"918E8B8A", x"88838080", x"7A7E7E79", x"787B7E7E",
									 -- x"7F7E7E7E", x"7F808284", x"817E7B7B", x"7B7A7B7D", x"83838486", x"898B8D8D", x"8F908F8F", x"92979998",
									 -- x"99999899", x"9DA09E9A", x"98949396", x"999B9D9F", x"9FA2A2A3", x"A7A8A9AC", x"AFB5BBBE", x"C0C1C1BF",
									 -- x"C3C5CACF", x"D0CDCBCB", x"CCCED0D2", x"D2D2D2D2", x"D2CFCCC9", x"C7C5C4C3", x"C0C0C2C5", x"CACED0D1",
									 -- x"D5D6D6D4", x"D2D2D2D1", x"CFCFCFCE", x"CED1D4D6", x"D3D7D9D9", x"D7D5D2CF", x"CAC9CBD0", x"D0CBC8C9",
									 -- x"C3C4C6C6", x"C5CACECB", x"CDD0CFCD", x"CDD0D0CD", x"CECDCDCE", x"D0D2D2D3", x"D4D5D7D6", x"D4D2D1D0",
									 -- x"CFCFCECB", x"C9C9C8C6", x"CBCBCAC9", x"C7C6C7C9", x"C3C3C3C3", x"C3C3C3C2", x"C2C3C4C5", x"C5C5C5C6",
									 -- x"C4C1C0C2", x"C4C3C0BC", x"BFC0C2C0", x"BEBDBFC1", x"BDBDBDBE", x"C2C7C5C1", x"C5C7CCD0", x"D1D0D1D4",
									 -- x"D4D4D5D5", x"D4D4D3D2", x"D5D7D8D6", x"D3D2D3D6", x"D7D8D9DA", x"DAD9D7D6", x"D8DADBDB", x"DADADADA",
									 -- x"DBDBDBDA", x"DADBDDDE", x"DCDCDDDD", x"DEDFE0E1", x"E1E0E0E1", x"E1E2E2E1", x"E2E2E3E2", x"E1DEDCDB",
									 -- x"D8D7D6D4", x"D2D1D0D0", x"CDCDCBC9", x"C6C4C5C6", x"C1BDBCBF", x"C0BCBABA", x"B6B5B2AE", x"AFB0AAA2",
									 -- x"A5A39F9C", x"9B9A9590", x"8E8E898D", x"8B8A8388", x"877E7C7F", x"7C787675", x"716F6F63", x"65626662",
									 -- x"5D5F5F5C", x"59575552", x"5252504D", x"4C4C4A46", x"4C44444B", x"4B464851", x"4A474443", x"474A4D4E",
									 -- x"4B4D4F50", x"4C4A4E55", x"51565553", x"585B5958", x"605D5D60", x"6262666D", x"6D6F6E6F", x"7171747B",
									 -- x"78808686", x"84878B8D", x"8A909697", x"97999B9C", x"97969498", x"9E9B9595", x"9E9A9A9B", x"98999D9E",
									 -- x"9E9D9893", x"97A0A29E", x"A09E9EA2", x"A5A5A5A6", x"AAAAABAA", x"A9AAAEB1", x"AAAEB0AF", x"AFB1AFAC",
									 -- x"AFADACAD", x"ACAAA9AB", x"A9A9ABAF", x"AEAAAAAE", x"AEA7A7A8", x"A4A6A7A1", x"A0A0A2A4", x"A4A1A0A2",
									 -- x"A5A4A3A1", x"A0A0A0A1", x"9E9A9B9C", x"9A98938B", x"9292908D", x"8A898A8B", x"89817C7E", x"7E7A7A7F",
									 -- x"77777471", x"7072716F", x"6D6A6767", x"66646364", x"615D595B", x"60615D57", x"55525356", x"56515052",
									 -- x"B2AFAAA6", x"A4A3A3A3", x"A1A0A0A0", x"A0A1A0A0", x"A19F9D9D", x"9D9E9D9D", x"9C9B9A9A", x"9A9B9B9B",
									 -- x"A2A3A6A7", x"A8A7A5A4", x"A1A2A29F", x"9B979798", x"96949290", x"8C878484", x"7D7C7A79", x"797A7E82",
									 -- x"81818180", x"80818384", x"827F7D7C", x"7C7B7B7C", x"80808285", x"898C8E8E", x"8D8F9091", x"95999B9A",
									 -- x"9B9B9B9C", x"9EA19F9B", x"98959497", x"9B9D9FA1", x"A2A5A5A6", x"AAACACB0", x"B9BCBFBF", x"C0C2C3C3",
									 -- x"C2C5CBD0", x"D1CECCCC", x"CDCECFD1", x"D2D2D2D2", x"D3D1CECA", x"C7C4C2C1", x"C1C3C5C7", x"C9CCCFD2",
									 -- x"D4D6D7D6", x"D5D5D4D2", x"CFD0D0CF", x"CFD0D2D3", x"D3D7DADA", x"D9D8D5D3", x"CFD2D4D4", x"D3D1CDCA",
									 -- x"C8C7C8C8", x"C7CBCECC", x"CDD2D5D3", x"D2D3D3D1", x"D1D0CFCF", x"D0D2D4D4", x"D6D7D8D8", x"D6D4D2D2",
									 -- x"D0D0CFCD", x"CCCCCCCA", x"CBCCCCCC", x"CAC9C9C9", x"C6C6C5C5", x"C5C5C4C4", x"C4C3C3C3", x"C4C5C5C5",
									 -- x"C1C0BFC1", x"C3C3C0BE", x"BDBFC0BF", x"BCBCBEC0", x"C0C0BFC0", x"C3C7C6C4", x"C7CCCFCE", x"CED0D1D0",
									 -- x"D4D3D3D3", x"D3D3D4D4", x"D4D4D4D3", x"D3D3D4D5", x"D4D6D8D8", x"D7D6D7D7", x"D9D9D9D9", x"D8D7D8D9",
									 -- x"DADADADA", x"D9DADBDC", x"DADADBDB", x"DCDDDEDE", x"DDDDDEDE", x"E0E0E1E1", x"E1E1E1E1", x"DFDDDBDA",
									 -- x"D8D8D7D5", x"D2CFCDCC", x"C9C9C9C7", x"C6C4C3C3", x"C3C1BFBF", x"BFBDBBBA", x"B5B1AEAF", x"B0AFABA7",
									 -- x"A2A1A09E", x"9D9A948E", x"8F918B8C", x"88888286", x"82828481", x"7B797976", x"71706F64", x"6460625E",
									 -- x"5F5F5D59", x"56565655", x"51514F4D", x"4D4E4C49", x"4846494F", x"4E47464B", x"49484849", x"4B4D4E4E",
									 -- x"494B4E50", x"4F4D4F52", x"53585654", x"585B5857", x"5B5B5E64", x"66656669", x"6A70706E", x"7175787C",
									 -- x"7C808484", x"84868A8C", x"8E939696", x"94939393", x"93939295", x"99979496", x"9997999C", x"9A9A9C9C",
									 -- x"9C9C9A98", x"9A9E9E9A", x"9D9FA2A4", x"A2A1A3A8", x"A7A8A8A7", x"A6A6A7A9", x"AAACAEAE", x"ADADABA8",
									 -- x"AAA9A8AA", x"AAA8A8AA", x"AAA8A8AB", x"A9A5A4A7", x"A4A2A2A3", x"A1A2A4A2", x"A1A0A0A2", x"A09E9E9F",
									 -- x"9E9D9B9B", x"9B9A9A9A", x"9B969595", x"9393928D", x"8B8C8B89", x"86858586", x"837F7D7F", x"7E7A7778",
									 -- x"73747370", x"6E6D6A67", x"6A676565", x"63615F60", x"5E5B5858", x"5B5C5955", x"55525356", x"55514F51",
									 -- x"B8B4AEAA", x"A8A8A7A6", x"A4A3A2A1", x"A2A2A2A2", x"A2A19F9D", x"9D9D9D9E", x"9C9C9B9A", x"9A9A9998",
									 -- x"A0A2A4A6", x"A7A6A5A4", x"9FA0A19F", x"9C9B9D9F", x"9D9C9A97", x"918B8787", x"847E7B7B", x"7B7A7E85",
									 -- x"80818281", x"7F7F8082", x"83807F80", x"80808081", x"84858688", x"8B8D8E8E", x"8E909294", x"989C9D9C",
									 -- x"9C9D9E9F", x"A0A1A09E", x"9A98979A", x"9DA0A2A3", x"A5A8A8A8", x"ADAEB0B4", x"BFC1C3C3", x"C3C5C5C5",
									 -- x"C2C6CCD2", x"D3D0CDCC", x"CDCDCED1", x"D3D4D3D2", x"D4D2CECB", x"C7C5C3C3", x"C3C5C8C8", x"C9CCD0D5",
									 -- x"D4D7D8D7", x"D6D5D3D1", x"D0D0D0D0", x"CFCFD0D1", x"D4D7DADB", x"DBDAD8D6", x"D4D9DCDA", x"D9DAD6D0",
									 -- x"CFCBCBCA", x"CACED1CF", x"CFD4D7D5", x"D3D4D5D4", x"D5D3D2D1", x"D2D3D5D5", x"D7D9DADA", x"D8D6D4D4",
									 -- x"D2D2D1CF", x"CECFCFCE", x"CCCDCECE", x"CDCBCAC9", x"C6C6C5C4", x"C4C3C3C4", x"C5C3C2C2", x"C3C4C5C4",
									 -- x"C3C2C2C3", x"C3C4C3C2", x"BEBFBFBE", x"BBBBBDBF", x"BFBFBFBF", x"C1C4C5C4", x"C4CBCECB", x"CCD2D4D1",
									 -- x"D4D3D3D2", x"D2D3D3D4", x"D3D2D0D0", x"D1D3D4D4", x"D2D5D7D7", x"D5D5D8DA", x"DAD9D8D6", x"D5D5D7D9",
									 -- x"D9DADAD9", x"D9D9D9DA", x"D9D9D9DA", x"DBDBDCDC", x"DCDCDDDD", x"DEDFDFDF", x"DFE0DFDF", x"DDDCDAD9",
									 -- x"D7D6D5D3", x"D0CDC9C8", x"C9C9C9C9", x"C9C7C5C3", x"C3C3C0BD", x"BDBDBAB8", x"B6B0ADB1", x"B2AFABAB",
									 -- x"A0A1A09F", x"9E9C9690", x"8E928B8A", x"85878082", x"7C81837D", x"787C7A71", x"70706E65", x"6460605C",
									 -- x"5E5E5B57", x"55555553", x"4E4C4A49", x"4A4C4A47", x"46474B4F", x"4D484546", x"46464748", x"494A4B4B",
									 -- x"48484A4D", x"4E4E4F50", x"52575553", x"57595858", x"5A5B6066", x"68676668", x"6770716C", x"70777A7B",
									 -- x"7E7E8083", x"85878A8D", x"8E929595", x"93939392", x"95969494", x"95939296", x"94929699", x"98979999",
									 -- x"9797989A", x"9C9D9D9D", x"9B9EA1A2", x"A09EA1A5", x"A4A5A6A5", x"A4A3A4A5", x"A6A6A7A9", x"A9A7A5A4",
									 -- x"A5A4A4A6", x"A6A5A5A6", x"A9A6A4A6", x"A5A19FA1", x"A0A2A19F", x"9F9E9DA0", x"A2A0A09F", x"9D9B9B9C",
									 -- x"9B9A9898", x"98989695", x"9490908F", x"8B8C8D8A", x"88898986", x"827F7E7E", x"7D7C7B7A", x"79777471",
									 -- x"6F70706E", x"6B6A6967", x"67646262", x"605D5B5B", x"5A595757", x"56565554", x"54525254", x"54504E50",
									 -- x"BAB6B0AD", x"ACACAAA7", x"A8A6A5A4", x"A3A3A3A2", x"A2A2A09E", x"9D9C9D9E", x"9D9C9C9B", x"9B9A9998",
									 -- x"9C9EA1A4", x"A5A5A4A3", x"A19E9B9B", x"9E9F9F9F", x"9F9F9E9A", x"938D8A89", x"8B847F7C", x"7A7A7E83",
									 -- x"7E808281", x"7E7D7E80", x"82818184", x"86878889", x"89888889", x"8B8D8D8E", x"92939596", x"999C9D9E",
									 -- x"9C9E9FA0", x"A1A1A2A2", x"9E9C9C9D", x"9FA1A3A4", x"A8ABABAB", x"B0B2B3B7", x"BDC0C4C7", x"C8C8C6C4",
									 -- x"C5C9CED2", x"D2D0CDCB", x"CCCCCDD1", x"D5D6D5D3", x"D1D0CECC", x"C9C8C7C7", x"C7C8CACB", x"CCCFD4D8",
									 -- x"D6D8D9D6", x"D4D3D1CE", x"CFCECECE", x"CECECFD1", x"D5D8DBDB", x"DBDAD9D7", x"D6DADEDF", x"E0E0DDD9",
									 -- x"D5D0CECD", x"CDD2D5D3", x"D4D6D6D4", x"D3D6D9D9", x"D8D6D4D4", x"D4D5D5D5", x"D8D9DADA", x"D9D8D6D5",
									 -- x"D4D4D2D0", x"CECFCFCE", x"CDCECECE", x"CDCBC9C8", x"C7C6C4C3", x"C2C2C3C3", x"C5C4C2C3", x"C4C5C4C3",
									 -- x"C5C6C6C4", x"C3C3C3C2", x"C0C0C0BE", x"BCBCBDBF", x"BEBFBFBF", x"C0C2C4C6", x"C3C7CACA", x"CCD1D3D3",
									 -- x"D3D3D3D2", x"D2D1D1D1", x"D2D0CFCE", x"CFD1D3D4", x"D3D5D6D7", x"D8D8DADC", x"D9D8D7D6", x"D5D6D7D9",
									 -- x"D9DADAD9", x"D9D8D8D9", x"D9DADADB", x"DBDBDBDB", x"DEDEDEDE", x"DEDDDEDE", x"DDDDDEDD", x"DCDBDAD9",
									 -- x"D6D5D4D2", x"D0CECBC9", x"CBCACACA", x"CAC9C6C4", x"C0C1BEBA", x"B9BBB9B6", x"B5B1AFB0", x"B1ADA8A6",
									 -- x"A2A19E9C", x"9B9B9996", x"8E928A89", x"8689807E", x"7D7B7A77", x"787E7A6D", x"6E6D6B65", x"6462625F",
									 -- x"5C5D5B58", x"5554514E", x"4C4A4746", x"48494743", x"48494A4B", x"4B4B4846", x"47474646", x"4647494B",
									 -- x"4B4A494A", x"4B4D5053", x"50555454", x"585B5B5C", x"5D5E6063", x"6566696B", x"6B72726F", x"7276787A",
									 -- x"7B7B7E83", x"86878B90", x"8D909292", x"92949595", x"94959392", x"94939295", x"95929497", x"95959999",
									 -- x"97959597", x"98989BA0", x"9B9B9B9D", x"9E9F9F9F", x"A1A1A2A2", x"A1A2A3A4", x"A3A1A2A6", x"A6A3A2A5",
									 -- x"A3A3A2A2", x"A1A0A0A0", x"A3A09E9F", x"9F9E9C9D", x"9DA19E9B", x"9E9B979B", x"9E9D9D9C", x"9A989797",
									 -- x"99979595", x"9594928F", x"8D8C8D8D", x"88868582", x"82838380", x"7D7A797A", x"78787572", x"7172716D",
									 -- x"6F6E6C68", x"65666769", x"64626160", x"5E5B5957", x"56575857", x"54535354", x"53515152", x"514E4D4E",
									 -- x"BAB7B3B1", x"B1AFACA9", x"ABA9A8A6", x"A5A4A3A2", x"A3A3A19F", x"9E9D9E9E", x"9E9D9D9C", x"9C9B9A99",
									 -- x"999B9EA1", x"A3A3A2A2", x"A4A19D9D", x"9FA1A1A0", x"9B9D9C99", x"94908E8E", x"8F8C857E", x"7C7E807F",
									 -- x"7F828382", x"807E7F81", x"82818387", x"8A8B8C8E", x"88878788", x"8A8C8E8F", x"95959697", x"999C9FA1",
									 -- x"A0A0A0A1", x"A0A0A1A3", x"A0A09FA0", x"A2A5A6A7", x"ACAFAEAF", x"B3B5B6BA", x"BCBFC4C9", x"CBC9C7C5",
									 -- x"C9CCD0D1", x"D0CECCCA", x"CACACCD1", x"D5D7D5D3", x"CFCFCECC", x"CBCACBCC", x"CDCDCDCE", x"D1D4D6D8",
									 -- x"D8D9D8D5", x"D2D1D0CE", x"CDCBCACB", x"CCCCCED2", x"D5D8DADB", x"DBDBDAD9", x"D7D8DDE3", x"E5E2E1E1",
									 -- x"DBD4D2D2", x"D1D4D7D5", x"D9D9D7D6", x"D8DBDCDB", x"D9D8D7D6", x"D6D6D5D4", x"D7D7D9DA", x"DAD9D7D6",
									 -- x"D4D4D3D0", x"CFD0D0CF", x"CFCFCECD", x"CCCAC9C8", x"C8C7C6C4", x"C3C3C3C4", x"C5C4C4C5", x"C6C6C5C3",
									 -- x"C4C6C6C3", x"C1C1C2C1", x"C1C1C1BF", x"BDBCBDBE", x"BFC0C1C1", x"C2C3C5C8", x"C7C5C7CB", x"CCCBCDD0",
									 -- x"D1D1D2D3", x"D3D1D0CF", x"D1D0CFCE", x"CDCFD1D3", x"D4D4D4D7", x"DADBDBDA", x"D7D7D6D7", x"D7D8D9D9",
									 -- x"DADADADA", x"D9D8D9D9", x"DADADBDB", x"DBDBDBDB", x"DDDEDEDE", x"DDDCDDDD", x"DCDCDCDC", x"DCDBDBDA",
									 -- x"D8D6D4D3", x"D1D0CECD", x"CBCAC8C7", x"C7C6C3C1", x"BDBEBDB9", x"B8BAB9B6", x"B1B1B0AE", x"ADABA59F",
									 -- x"A3A19E9A", x"98999895", x"8F918989", x"898D827E", x"827B7878", x"797A7770", x"6B6A6664", x"62636261",
									 -- x"5B5B5956", x"5453504C", x"4D4C4A48", x"494B4945", x"49494949", x"4C4F4D47", x"4A4A4A49", x"494A4B4D",
									 -- x"4C4D4D4C", x"4C4E5254", x"50555556", x"5B5D5D60", x"5F606161", x"63676B6D", x"70737374", x"7675767B",
									 -- x"777A8084", x"86888C91", x"8F90908E", x"8F919292", x"8F908F8F", x"93949293", x"95939598", x"96959898",
									 -- x"99959495", x"9493959B", x"999A9A9B", x"9C9D9E9D", x"9E9E9D9D", x"9D9FA1A3", x"A4A1A0A3", x"A3A1A2A5",
									 -- x"A1A1A09F", x"9E9D9D9C", x"9C999898", x"99999999", x"979A9696", x"9B9A9597", x"96979897", x"95939291",
									 -- x"918F8E8E", x"8E8D8B89", x"8A898B8B", x"8683827F", x"7A7B7B7A", x"78787979", x"7374716D", x"6D6F6E6B",
									 -- x"706D6863", x"605F6062", x"61605F5E", x"5D5B5855", x"51535655", x"53505052", x"51504F4F", x"4E4C4B4B",
									 -- x"BAB8B5B4", x"B4B2AFAD", x"ADACAAA9", x"A7A6A4A3", x"A4A4A3A1", x"A0A09F9F", x"9F9E9D9D", x"9D9C9B9B",
									 -- x"9B9DA0A3", x"A4A4A3A2", x"A1A2A2A0", x"9D9C9FA1", x"97999997", x"95959594", x"96958E87", x"85888782",
									 -- x"82838483", x"81808081", x"84838487", x"8A8B8C8D", x"8D8C8A8A", x"8B8D8E8E", x"93939597", x"9A9CA0A4",
									 -- x"A4A3A2A2", x"A1A0A0A2", x"A0A2A3A3", x"A5A9ACAC", x"ADB1B1B1", x"B4B5B5B9", x"C0C1C4C9", x"CBCAC9C8",
									 -- x"CACDD0D0", x"CFCDCBC9", x"C7C8CACD", x"D1D3D2D2", x"CECECECD", x"CBCBCCCE", x"D2D2D2D3", x"D5D6D6D6",
									 -- x"D7D9D8D4", x"D2D1D0CF", x"CAC8C7C9", x"C9C9CCD0", x"D2D5D8D9", x"D9DBDBDA", x"D8D7DBE2", x"E4E1E0E2",
									 -- x"DED8D6D6", x"D4D6D8D7", x"D9D8D8DA", x"DDDEDBD8", x"DAD9D9D8", x"D8D7D5D4", x"D6D6D7D9", x"D9D9D7D5",
									 -- x"D3D3D2CF", x"CFD0D1D0", x"D1CFCECC", x"CCCBC9C8", x"C7C6C5C4", x"C3C3C3C3", x"C5C6C7C8", x"C8C8C6C6",
									 -- x"C6C8C7C4", x"C3C4C4C2", x"C0C0C0BF", x"BEBDBDBE", x"BFBFC0C1", x"C2C2C4C6", x"C6C2C3C9", x"CBC9CACF",
									 -- x"CDCED0D2", x"D3D2D1D0", x"D0CFCECD", x"CCCDCFD2", x"D2D1D1D4", x"D8DAD8D6", x"D5D5D5D7", x"D8D9DADA",
									 -- x"DADADADA", x"D9D9D9DA", x"DADADBDB", x"DBDADAD9", x"DADBDCDC", x"DBDADBDD", x"DBDBDBDB", x"DBDBDBDA",
									 -- x"D8D6D3D1", x"D0CFCDCB", x"CCCAC8C6", x"C5C3C2C1", x"BEBEBDBB", x"BABABAB9", x"B0B3B2AF", x"AEADA8A0",
									 -- x"A2A2A09C", x"99979390", x"8D8E8688", x"898B817E", x"837C7B7B", x"75717273", x"6B696464", x"60636161",
									 -- x"5B5A5754", x"5354524F", x"4D4D4C4B", x"4B4C4A47", x"45464648", x"4C4F4B45", x"4848494A", x"4B4B4A4A",
									 -- x"4A4C4E4E", x"4D4E4F4F", x"4F535556", x"5A5B5A5D", x"5D606262", x"64696C6C", x"6F727274", x"7674747A",
									 -- x"777D8385", x"86898C8E", x"90908F8E", x"8F929291", x"9092908F", x"92938F8F", x"908F9498", x"96949391",
									 -- x"92919294", x"94929395", x"94999E9C", x"99999DA0", x"9E9D9C9B", x"9C9D9FA0", x"A09E9D9D", x"9D9C9D9F",
									 -- x"9D9E9D9C", x"9B9B9B9A", x"99979696", x"96969696", x"95969494", x"97969290", x"91939493", x"91908F8D",
									 -- x"8B8B8B8A", x"89898989", x"87858686", x"82818280", x"7C7B7978", x"77777675", x"6E6F6F6D", x"6D6E6B67",
									 -- x"6A676463", x"615F5E5E", x"5D5D5D5B", x"5A595754", x"4D505252", x"504E4D4E", x"4D4D4D4C", x"4B4A4949",
									 -- x"B8B7B6B5", x"B4B3B2B1", x"AEADACAB", x"AAA8A6A4", x"A6A5A4A4", x"A4A3A2A0", x"A09F9E9D", x"9D9C9C9B",
									 -- x"9C9DA0A3", x"A4A4A4A3", x"9FA0A19F", x"9C9B9D9F", x"999A9A98", x"999B9C9B", x"9F9B9692", x"918F8B87",
									 -- x"86868685", x"83828282", x"88868688", x"8A8A8A8C", x"9391908F", x"8F8E8D8C", x"91919498", x"9B9DA1A5",
									 -- x"A5A4A4A5", x"A5A3A2A3", x"A2A5A6A7", x"A9ADB0B0", x"B1B5B5B5", x"B8B7B6B9", x"C1C1C4C9", x"CCCBCACA",
									 -- x"C8CCCFCF", x"CFCECBC8", x"C5C6C6C7", x"C9CBCDCF", x"CBCCCDCC", x"CACACCCE", x"D3D4D6D7", x"D7D7D6D5",
									 -- x"D6D8D7D4", x"D1D0CECC", x"C9C6C6C8", x"C8C6C8CD", x"CED1D3D4", x"D5D6D7D6", x"D4D5D9DC", x"DEDEDDDD",
									 -- x"DDD8D9DA", x"D7D7DADA", x"D9D9DADC", x"DDDDDBD9", x"DCDBDAD9", x"D8D8D6D5", x"D7D7D7D8", x"D9D8D6D4",
									 -- x"D2D2D0CD", x"CDCECFCE", x"CFCDCCCB", x"CBCAC9C8", x"C5C5C4C4", x"C3C3C2C2", x"C6C8CACA", x"C9C8C9CA",
									 -- x"CACCCBC7", x"C6C7C6C3", x"BFBFC0C0", x"C0C0C0C0", x"BFBEBEC0", x"C1C0C0C2", x"C3C1C2C6", x"C9C8C9CB",
									 -- x"CCCDCFD1", x"D2D2D2D1", x"CFCDCBCA", x"CBCDCECF", x"D0CFCFD1", x"D3D5D5D4", x"D4D3D3D5", x"D7D9D9D9",
									 -- x"DADADAD9", x"D8D8DADB", x"DADADBDB", x"DBDAD9D9", x"D9DADBDB", x"D9D9DADB", x"DBDBDBDA", x"DADAD9D9",
									 -- x"D7D5D2D1", x"D0CFCCCA", x"CCCCCBC8", x"C6C4C3C2", x"C1C0BFBF", x"BDBAB9BA", x"B3B3B2B1", x"B0ADA9A5",
									 -- x"A3A3A29E", x"9B989490", x"8D8C8588", x"87877F81", x"817B7A7A", x"726D6F71", x"6C6A6467", x"62656060",
									 -- x"5B5A5856", x"56565450", x"4C4E4E4C", x"4B4A4947", x"43444647", x"4A4A4845", x"45454647", x"4A4B4A4A",
									 -- x"4A4C4D4D", x"4F50504D", x"4E535456", x"5A59595C", x"5A5F6363", x"666C6E6C", x"6F747574", x"75757578",
									 -- x"79808484", x"868B8D8A", x"8E8E8F8F", x"92949391", x"9094928F", x"90908D8D", x"8D8D9297", x"9491908E",
									 -- x"8C8C8E91", x"92939393", x"91979C9A", x"97979B9F", x"9D9C9B9B", x"9B9C9D9E", x"9A9B9A99", x"98999A99",
									 -- x"999A9A98", x"97999896", x"95959594", x"92929293", x"94929394", x"92918F8B", x"8D8F908E", x"8C8D8C8A",
									 -- x"88898987", x"85848586", x"807D7E7E", x"7B7C7E7D", x"7C797676", x"7675716E", x"6B6B6C6C", x"6C6B6764",
									 -- x"635F5E61", x"62615E5D", x"58595856", x"56575552", x"4E4E4E4E", x"4D4C4C4B", x"4A4A4A49", x"48484747",
									 -- x"B7B6B5B4", x"B3B3B3B3", x"AEAEAEAD", x"ACABA8A6", x"A8A6A5A5", x"A6A6A4A1", x"A1A09E9C", x"9C9C9B9B",
									 -- x"97999DA0", x"A2A3A2A2", x"A19F9D9D", x"9F9F9D9B", x"9D9D9C9B", x"9C9F9F9E", x"A39C9898", x"968F8987",
									 -- x"8C8B8A88", x"87868584", x"8B89888A", x"8B8A8B8C", x"90909090", x"908F8E8C", x"90909499", x"9B9CA0A4",
									 -- x"A4A3A4A8", x"A9A7A5A5", x"A5A8A9A9", x"ABAFB1B1", x"B7BBBBBB", x"BDBCBABD", x"BEBFC3CA", x"CECDCBCA",
									 -- x"C5CACECF", x"CFCFCCC8", x"C5C4C3C3", x"C3C6C9CC", x"C8CACBCA", x"CACACDCF", x"D1D5D8D9", x"D8D6D6D7",
									 -- x"D5D7D7D4", x"D0CDCAC8", x"C9C6C6C8", x"C7C4C5C9", x"CBCED0D0", x"D0D1D1D0", x"CFD3D6D6", x"D8DCDBD8",
									 -- x"DAD7D9DB", x"D9D9DCDD", x"DDDCDDDD", x"DDDCDDDE", x"DEDCDAD9", x"D9D8D8D7", x"D8D7D7D8", x"D8D7D5D2",
									 -- x"D2D1CFCB", x"CACBCBCA", x"CBCACACA", x"CACAC8C7", x"C6C6C6C6", x"C6C5C4C4", x"C7C9CBCB", x"C9C9CBCD",
									 -- x"CCCDCBC7", x"C6C7C4C0", x"BFC0C1C2", x"C3C3C3C2", x"C2C0BFC2", x"C3C1C0C1", x"C4C5C5C4", x"C5C6C5C3",
									 -- x"CDCECFD0", x"D1D1D1D1", x"CECBC8C9", x"CBCECDCC", x"CFCFCFCF", x"D0D2D3D5", x"D3D2D2D3", x"D5D7D8D8",
									 -- x"DAD9D9D8", x"D7D8DADB", x"DBDBDCDC", x"DCDBDAD9", x"DADBDCDB", x"D9D8D9DA", x"DBDBDBDA", x"D9D8D8D8",
									 -- x"D7D6D4D4", x"D4D2CFCC", x"CBCCCCC9", x"C6C3C3C3", x"C4C1C1C2", x"BFBAB8BA", x"B4B0AEB0", x"AEA9A6A6",
									 -- x"A5A5A39F", x"9C9A9795", x"908F888B", x"87878187", x"817A7777", x"7472716E", x"6D6C666A", x"65686162",
									 -- x"5A5B5A5A", x"5958534E", x"4E50514F", x"4B494745", x"47484949", x"4948494B", x"4A484647", x"4B4E5050",
									 -- x"504F4D4D", x"51555450", x"50545759", x"5D5C5B5F", x"595F6263", x"666D706E", x"727A7B76", x"777A7979",
									 -- x"7A818482", x"868E8F89", x"8D8E8F8F", x"91918E8A", x"898F8E8B", x"8C8D8E91", x"918F9396", x"93929392",
									 -- x"8D8D8D8D", x"8F91918F", x"91949695", x"96999A9A", x"99989899", x"9A9A9A9A", x"979A9B99", x"999B9B98",
									 -- x"97999896", x"95969593", x"8E90908F", x"8D8D8D8E", x"8B898F91", x"8D8D8F8B", x"888A8A87", x"86878785",
									 -- x"83848481", x"7D7B7C7F", x"7A777879", x"77787875", x"73716F70", x"73736F6B", x"6B696869", x"69676462",
									 -- x"615C5A5C", x"5E5C5A58", x"54555553", x"53545350", x"514F4D4C", x"4C4C4B4B", x"48494847", x"47474646",
									 -- x"B9B7B6B6", x"B6B5B2B0", x"B2B1AFAC", x"ABABAAA8", x"A8A7A7A7", x"A8A7A5A4", x"A2A09E9D", x"9B99999A",
									 -- x"969A9C9D", x"A0A3A29E", x"A29F9D9E", x"9F9F9FA0", x"969DA1A1", x"9F9FA0A0", x"9DA2A29E", x"9A97928D",
									 -- x"8F8E8F8F", x"8D8A8A8C", x"8F91918D", x"8A8A8C8C", x"91949796", x"94928F8D", x"91939597", x"999CA1A5",
									 -- x"A4A6A8A7", x"A8A8A7A6", x"AAA7AAB0", x"B1AEB0B7", x"BCBCBCBD", x"BDBEBEBF", x"C2C4C7CA", x"CCCCCBCA",
									 -- x"C4C7CACB", x"CCCDCAC7", x"C4C3C4C5", x"C5C2C2C3", x"C4C5C6C8", x"C8C7C6C5", x"CCD3D9DA", x"D8D6D5D3",
									 -- x"D4D2D1D1", x"D0CDCAC9", x"C4C3C2C3", x"C2C1C3C6", x"C5C6C9CE", x"CECBC9C8", x"C9CCD2D7", x"D7D5D4D7",
									 -- x"D3D7DBDB", x"D9D8DBDF", x"DEDDDDDE", x"DFDEDBD9", x"DBDBDAD9", x"D8D8D7D4", x"D4D5D6D6", x"D5D4D3D2",
									 -- x"D2CDC9C9", x"C9C9C9CB", x"CBCAC8C8", x"C8C8C8C7", x"C6C6C7C8", x"C7C4C5C8", x"C9CACCCD", x"CDCECFD0",
									 -- x"CFCECCCA", x"C9C8C4C0", x"C2C1C1C2", x"C4C5C4C3", x"C1C1C1C2", x"C1C1C1C1", x"C4C4C4C3", x"C3C3C5C7",
									 -- x"CBCCCECE", x"CDCDCFD0", x"CECFCCC8", x"C7CCCFCF", x"CCCECFCE", x"CFD1D3D2", x"D6D4D2D1", x"D2D4D5D6",
									 -- x"D6D8DADA", x"DAD9DADB", x"DCDDDEDC", x"DBDCDCDB", x"DDDADBDE", x"DBD9DADA", x"DEDCDAD9", x"D9D9D7D6",
									 -- x"D6D7D7D3", x"CFCFD0D1", x"CAC9C8C7", x"C6C4C3C2", x"C6C1BEBE", x"BDB9B9BB", x"BAB6B1AF", x"AFACA8A5",
									 -- x"A4A2A19D", x"999A9992", x"8F8E8B88", x"85838282", x"837E7975", x"74726E6B", x"6C6B6865", x"65635F5A",
									 -- x"5D5C5A59", x"58575451", x"52535350", x"4B484A4D", x"48484847", x"4747494A", x"47474848", x"484A4B4D",
									 -- x"4E4D4D4F", x"50515457", x"52575F5F", x"5A60645F", x"62646667", x"696D7174", x"72747677", x"7676787A",
									 -- x"7C7D8085", x"898A8A8B", x"8D8D8C8C", x"8D8F8E8B", x"8C8F8C88", x"8A8F8F8B", x"908D8C8E", x"9193928F",
									 -- x"8E8F8D8B", x"8C909394", x"928D9297", x"92919697", x"90949797", x"97979796", x"95979796", x"95959799",
									 -- x"95949494", x"94939392", x"908D8F90", x"8D8D8B86", x"8A8A8B8C", x"8B89888A", x"86878582", x"82848482",
									 -- x"827F7C7A", x"7B7B7B7A", x"7C7B7876", x"73727171", x"726E6C6E", x"706E6B69", x"69686562", x"5F5F6163",
									 -- x"5E5C5B5B", x"5B595858", x"53545453", x"52515152", x"4C4D4C49", x"4A4E4F4D", x"48484746", x"44434344",
									 -- x"BBB9B6B6", x"B6B6B4B3", x"B1B1AFAD", x"ADAEAEAC", x"A9A9A9AA", x"AAA9A7A5", x"A5A3A09E", x"9C999898",
									 -- x"97999B9D", x"A0A2A19F", x"A19F9EA0", x"A09E9C9C", x"9A9EA1A0", x"9FA0A2A2", x"A2A4A4A1", x"A0A09C97",
									 -- x"9A938E8F", x"91908C8A", x"8F919290", x"8E8F8F8E", x"91949797", x"96969594", x"92949697", x"999B9FA1",
									 -- x"A1A6AAAA", x"A9AAACAD", x"AAA9AAAE", x"AFAFB2B7", x"BEBEBEBF", x"BFC0C0C1", x"C1C4C8CB", x"CBCBC9C9",
									 -- x"C1C3C4C5", x"C6C7C6C3", x"C2C1C1C3", x"C2C0BFC0", x"BEBEBFBF", x"C0C0C0C1", x"C6CCD3D5", x"D6D7D7D6",
									 -- x"D4D3D2D1", x"D1CECAC7", x"C3C2C2C1", x"C0BFC1C3", x"C2C3C5C9", x"C9C7C5C5", x"C5C8CED3", x"D4D1CFCF",
									 -- x"D0D2D5D7", x"D8D8D9D9", x"DBDBDCDB", x"DAD9D9D8", x"DBDBD9D7", x"D6D6D5D3", x"D2D2D2D2", x"D1D0CFCF",
									 -- x"CFCDCBCA", x"C8C7C9CB", x"C8C7C7C7", x"C7C7C6C5", x"C6C6C7C8", x"C7C6C7C9", x"C9CBCCCD", x"CDCECECF",
									 -- x"CECFCECC", x"CAC9C6C3", x"C4C3C2C2", x"C3C4C4C3", x"C1C1C2C2", x"C2C2C2C2", x"C2C3C4C4", x"C4C5C7C8",
									 -- x"CBCBCBCC", x"CDCECECE", x"CAC9C7C6", x"C7CBCCCB", x"CCCECECD", x"CED0D2D2", x"D1D1D2D3", x"D5D6D6D6",
									 -- x"D6D6D7D8", x"D9DADADA", x"D7DBDDDC", x"DADADBDB", x"DCD8DADD", x"DBDADBDA", x"DBDAD9D9", x"D8D7D6D5",
									 -- x"D6D7D6D3", x"D1D1D0CF", x"CBC9C7C5", x"C3C3C4C5", x"C2C0BEBD", x"BBBABABC", x"B6B3B0AF", x"AEABA6A3",
									 -- x"A5A2A19F", x"9B9A9791", x"8F8D8B89", x"86838180", x"817D7874", x"716E6B69", x"68696865", x"63615E5B",
									 -- x"5C5A5857", x"56565554", x"5252514F", x"4C4B4C4D", x"4B474446", x"4A4C4A47", x"4C4B4A48", x"48494C4E",
									 -- x"50505051", x"50505153", x"54585D5E", x"5D61625F", x"61636668", x"6A6C6F71", x"70727576", x"7676787A",
									 -- x"7E7F8081", x"83858483", x"898A8A8A", x"8C8E8D8A", x"8D8C8B8A", x"8A8B8B8C", x"8E8D8B8C", x"8E8F8D8B",
									 -- x"8C8D8C8B", x"8D909291", x"948E9195", x"91909393", x"8F929594", x"93939392", x"8F909191", x"90909090",
									 -- x"9391908F", x"8F908E8D", x"8B888A8B", x"8A8A8A86", x"85848386", x"87878687", x"8384837F", x"7E7E7E7D",
									 -- x"7D7C7B7A", x"78777777", x"74737271", x"7170706F", x"706C696B", x"6B696563", x"65636262", x"62626160",
									 -- x"5C5A5A5B", x"5A585757", x"50515150", x"4F4F4F50", x"4C4E4E4C", x"49484746", x"47474544", x"43434343",
									 -- x"BCB9B6B5", x"B5B6B6B5", x"B1B1B0AF", x"AFB1B0AF", x"ABABACAD", x"ADABA9A8", x"A8A5A3A1", x"9E9B999A",
									 -- x"9998989C", x"9F9F9FA0", x"A19F9E9F", x"9F9C9A9A", x"9E9F9F9D", x"9DA0A2A3", x"A4A5A4A3", x"A6A9A7A3",
									 -- x"A49D9694", x"9493908E", x"8E919293", x"94949492", x"91939595", x"96989999", x"93939496", x"989A9D9E",
									 -- x"9FA6ABAB", x"AAACAFB2", x"AEAFAFAF", x"B0B4B8BC", x"BFC0C0C0", x"C1C2C2C2", x"C2C6CACD", x"CECDCBCA",
									 -- x"C3C3C3C2", x"C3C4C5C4", x"C0C0C0C1", x"C1BFBEBE", x"BCBBBABA", x"BABCBFC0", x"C1C6CBCF", x"D3D5D6D5",
									 -- x"D2D2D2D1", x"D0CDC9C5", x"C3C1C0C0", x"BEBCBDC0", x"C1C1C2C4", x"C5C4C3C4", x"C4C5C9CD", x"D0CFCDCD",
									 -- x"CCCDCFD3", x"D7D8D6D4", x"D7D8D9D8", x"D6D5D7D9", x"DCDCDAD7", x"D6D7D6D4", x"D1D1D0CF", x"CECECDCC",
									 -- x"CBCAC9C8", x"C6C4C6C9", x"C5C4C4C5", x"C6C6C5C4", x"C6C6C8C9", x"C9C8C9CB", x"CBCCCECE", x"CECFCFD0",
									 -- x"CDD0D1CE", x"CCCAC8C6", x"C6C4C3C2", x"C3C4C4C3", x"C2C2C2C2", x"C2C2C3C3", x"C0C1C3C4", x"C4C5C6C7",
									 -- x"CAC9C8C9", x"CBCCCBC9", x"CAC6C5C7", x"CACAC9C9", x"CBCCCCCC", x"CCCFD1D1", x"D0D0D1D3", x"D5D7D7D7",
									 -- x"D6D4D4D5", x"D8DAD9D8", x"D3D8DCDB", x"D9D9DADB", x"DCD8D9DC", x"DBDBDCD9", x"D9D9DAD9", x"D8D7D7D6",
									 -- x"D6D7D6D4", x"D3D2D0CE", x"CDCCC9C6", x"C4C3C2C2", x"BEBEBDBB", x"B9BABBBB", x"B2B2B1AF", x"ADAAA6A3",
									 -- x"A6A1A1A1", x"9C989590", x"8E8D8C8A", x"8784807E", x"7E7C7875", x"716E6D6C", x"66686966", x"63615F5D",
									 -- x"5C5A5856", x"55555555", x"52514F4E", x"4D4D4C4B", x"4D494648", x"4C4F4D4A", x"4C4B4948", x"494C5154",
									 -- x"50505153", x"53525355", x"595B5C5E", x"63636060", x"6264686A", x"6B6C6D6E", x"72747677", x"77797B7D",
									 -- x"7D80807F", x"80848483", x"8587888A", x"8C8E8D8A", x"8C8A898A", x"8886878A", x"8A8A8A8B", x"8B8A8988",
									 -- x"8A8B8B8C", x"8E90908F", x"928C8D90", x"8F8F908E", x"8F919291", x"8F8F8E8D", x"8D8E8F90", x"8F8F8E8D",
									 -- x"8F8C8A89", x"8B8B8987", x"88858788", x"87888885", x"85817F80", x"82817F7F", x"7E7F7E7B", x"7A7A7A7A",
									 -- x"76787877", x"75737272", x"706E6D6E", x"70706F6D", x"6C686667", x"69686564", x"5F5D5E61", x"6565605C",
									 -- x"5B5A5A5A", x"58555455", x"5050504F", x"4E4E4F50", x"494A4A4A", x"47444446", x"46444241", x"41414140",
									 -- x"BBB9B6B4", x"B4B4B4B4", x"B3B3B2B1", x"B1B2B1AF", x"AEAEAEAE", x"AEADACAB", x"A7A5A4A3", x"A19F9E9F",
									 -- x"9D9A999D", x"9F9E9FA1", x"A29F9D9D", x"9C9B9B9D", x"A09E9C9B", x"9B9D9E9F", x"A2A3A3A4", x"A7ABABA8",
									 -- x"A8A7A49E", x"98939394", x"8F909294", x"96979795", x"95969696", x"97999B9A", x"94939294", x"969A9C9D",
									 -- x"9FA5AAAA", x"AAACAFB2", x"B2B4B4B1", x"B2B7BCBE", x"C0C0C0C1", x"C2C2C2C2", x"C4C6C9CE", x"D1D0CDCA",
									 -- x"C6C5C3C2", x"C2C3C4C4", x"C0C0C0C1", x"C1BFBEBD", x"BCBAB9B8", x"BABCBFC1", x"C2C4C8CB", x"CED0D0D0",
									 -- x"D2D1D0CF", x"CECCC9C5", x"C3C1BFBE", x"BCBBBBBD", x"BFBFBFC0", x"C1C1C2C3", x"C4C3C3C5", x"C9CCCCCC",
									 -- x"C8C8CACE", x"D2D4D3D1", x"D3D4D5D4", x"D4D4D6D7", x"D8D9D9D7", x"D7D7D5D2", x"CECECECE", x"CDCCCBCA",
									 -- x"C6C5C5C5", x"C3C2C3C5", x"C2C2C3C4", x"C5C5C4C3", x"C6C8CACB", x"CBCACBCD", x"CFD0D1D1", x"D1D1D1D2",
									 -- x"CFD1D1CF", x"CDCCC9C7", x"C7C5C3C3", x"C3C4C4C4", x"C2C2C2C2", x"C2C3C4C4", x"C0C1C2C3", x"C4C4C4C4",
									 -- x"C8C8C7C8", x"C9C9C8C6", x"CAC7C6C9", x"CAC8C6C8", x"C8C9C9C9", x"CACCCFD1", x"D2D1D0D0", x"D2D4D6D7",
									 -- x"D5D4D4D4", x"D6D8D8D8", x"D3D7DBDA", x"DADADBDB", x"DCD9D9DB", x"DADBDBD8", x"D9DADCDC", x"DAD9D9D9",
									 -- x"D8D7D5D4", x"D4D4D1CD", x"CBCBCAC9", x"C7C5C3C1", x"BCBDBCB9", x"B9BBB9B5", x"B1B3B3B0", x"ADAAA8A5",
									 -- x"A6A0A0A1", x"9C979491", x"908E8C8A", x"8784807D", x"79797875", x"72707070", x"6A6B6A67", x"64636260",
									 -- x"5D5C5A58", x"56555453", x"5251504F", x"4D4B4A49", x"4B4B4B4A", x"4A4C4D4F", x"4A494949", x"4B4E5356",
									 -- x"51515255", x"55555759", x"5F605C5F", x"68666061", x"64666A6C", x"6C6D6E70", x"73747677", x"78797C7D",
									 -- x"7B7F817F", x"7F838583", x"82858788", x"8B8C8B88", x"8A898787", x"86858586", x"85868889", x"8A898989",
									 -- x"8988888A", x"8D8F8E8D", x"8C89888B", x"8B8B8C8C", x"8E8F8F8D", x"8C8C8B8A", x"8B8D8F8F", x"8D8C8C8C",
									 -- x"8A878585", x"88888582", x"87838484", x"82838480", x"827F7E7F", x"7F7D7A7A", x"78777675", x"76777675",
									 -- x"73747473", x"72706E6D", x"6E6D6C6D", x"6F6E6B68", x"6A666363", x"64656463", x"5A5A5C60", x"64635E59",
									 -- x"5B5B5A5A", x"56525151", x"5151504F", x"4E4E4E4F", x"4B474445", x"44424449", x"45423F3F", x"40403E3C",
									 -- x"BBBAB8B6", x"B5B5B4B4", x"B4B4B4B2", x"B2B3B2B0", x"B0B0B0B0", x"AFAFAFAF", x"A7A5A4A5", x"A4A2A1A3",
									 -- x"A29E9D9F", x"A19F9FA1", x"A09E9D9D", x"9C9C9D9F", x"A19E9C9B", x"9C9C9B9B", x"9FA2A4A5", x"A7A9A9A9",
									 -- x"A8ABACA6", x"9C959496", x"91919294", x"96979797", x"999A9998", x"999C9D9D", x"97959393", x"95989B9C",
									 -- x"A1A5A7A9", x"ABAEB0B0", x"B3B5B5B1", x"B1B6BBBB", x"C0C0C1C2", x"C2C3C3C3", x"C3C3C5CA", x"D0D1CDC9",
									 -- x"C5C3C0BF", x"BFC0C0C1", x"C1C1C1C1", x"C1C0BEBC", x"B9B8B7B7", x"B8BABCBE", x"C2C3C5C8", x"CACBCCCC",
									 -- x"D1D1D0CD", x"CDCDCBC7", x"C3C0BEBD", x"BCBABABB", x"BBBBBBBB", x"BCBEC0C1", x"C2C0BEBF", x"C3C6C7C6",
									 -- x"C3C4C5C8", x"CACDCECE", x"CFCFD0D1", x"D2D2D1CF", x"D0D2D4D4", x"D4D4D2CE", x"C9C9CACA", x"CAC9C7C6",
									 -- x"C4C2C0C1", x"C2C1C1C1", x"C0C1C3C4", x"C4C4C4C4", x"C7C9CBCC", x"CCCCCDCE", x"D0D1D2D2", x"D2D2D3D3",
									 -- x"D2D2D1CF", x"CECDC9C5", x"C8C6C3C3", x"C4C4C4C4", x"C3C3C3C3", x"C3C3C4C4", x"C0C0C1C2", x"C3C4C4C4",
									 -- x"C4C5C7C7", x"C7C6C6C7", x"C7C5C5C7", x"C5C2C3C6", x"C5C5C5C6", x"C8CACDD0", x"D1D0CFCF", x"D1D3D4D5",
									 -- x"D5D5D6D5", x"D5D5D6D8", x"D7D9D9D9", x"DADCDCDA", x"DCD9DADB", x"DADBDCD8", x"DADBDDDD", x"DCDBDBDB",
									 -- x"DAD8D6D4", x"D4D5D3CF", x"C8C8C8C8", x"C7C6C5C4", x"BEBEBCBA", x"BBBCB7B1", x"B2B4B3AF", x"ABAAA9A7",
									 -- x"A69F9EA0", x"9B979593", x"928F8C89", x"8784817F", x"78797875", x"716E6E6F", x"6D6B6865", x"64646360",
									 -- x"5C5C5D5C", x"5A575553", x"53535352", x"4E4C4B4B", x"4B4B4A49", x"494A4D4E", x"4C4C4D4E", x"4E4F5152",
									 -- x"54535354", x"55555759", x"62625D5F", x"68676062", x"6567696B", x"6C6D7072", x"73737373", x"7476787A",
									 -- x"7A7E807F", x"7E808180", x"81838586", x"87898885", x"898A8784", x"85898782", x"82848789", x"89898A8B",
									 -- x"88868688", x"8A8B8C8C", x"88888787", x"8888888B", x"8B8B8A88", x"87888887", x"85878988", x"85848587",
									 -- x"85838183", x"8686827F", x"827E7E7E", x"7C7D7D7A", x"7A7A7B7D", x"7C7A7879", x"76727070", x"72726F6D",
									 -- x"72706E6E", x"6F6F6C69", x"6C6A696A", x"6C6B6763", x"6B686360", x"5F5F5F5D", x"5A5B5D5F", x"605E5A57",
									 -- x"5B5A5958", x"55514F50", x"5150504E", x"4C4B4C4C", x"51494242", x"43424244", x"45423F3F", x"3F3F3D3B",
									 -- x"BBBABAB8", x"B7B6B5B5", x"B4B5B5B4", x"B5B7B6B4", x"B3B4B4B3", x"B2B2B2B3", x"AAA8A8A8", x"A7A4A3A4",
									 -- x"A3A19E9F", x"9F9F9E9F", x"9F9E9FA1", x"A09E9D9E", x"A09E9D9E", x"9E9C9C9C", x"A0A3A6A8", x"A8A9A9AA",
									 -- x"ABACABA6", x"A19C9894", x"95949495", x"95959597", x"98999998", x"9A9E9F9E", x"9C9A9795", x"95979A9D",
									 -- x"A3A4A6A8", x"ADB2B3B1", x"B3B6B6B3", x"B3B6B9BA", x"C0C1C2C3", x"C3C3C3C3", x"C3C2C3C8", x"CED1CECA",
									 -- x"C5C1BFBE", x"BDBDBDBE", x"C0C1C0C0", x"C0C0BDBA", x"B7B7B7B7", x"B7B8BABB", x"BEBFC2C5", x"C7C8C9CC",
									 -- x"D0D0CFCC", x"CCCECDC9", x"C3C0BDBC", x"BBB9B8B9", x"B9BABAB9", x"BABDBFBF", x"BDBEBDBE", x"C0C2C1BE",
									 -- x"C1C1C2C3", x"C5C7CACC", x"CBCACBCC", x"CDCCC9C6", x"C9CCD0D1", x"D2D2CFCC", x"C6C6C7C7", x"C7C6C5C4",
									 -- x"C3C0BEBF", x"C1C1C0C0", x"C0C1C3C3", x"C3C3C4C4", x"C6C9CCCC", x"CCCDCECD", x"D0D1D2D2", x"D2D2D3D3",
									 -- x"D5D3D1CE", x"CECEC9C5", x"C8C6C4C3", x"C4C4C4C3", x"C3C3C3C3", x"C3C3C3C3", x"C0C0C0C1", x"C3C4C5C5",
									 -- x"C1C3C6C6", x"C6C5C6C7", x"C3C3C4C4", x"C2C1C3C6", x"C3C2C3C5", x"C7C8CBCE", x"CCCDCED1", x"D3D4D3D3",
									 -- x"D4D6D7D6", x"D4D4D5D7", x"DAD9D9D9", x"DBDDDDDA", x"D9D8DBDB", x"DADCDEDB", x"DBDCDDDD", x"DCDCDCDC",
									 -- x"DBDAD7D5", x"D5D6D4D0", x"CDCBC8C4", x"C2C2C2C3", x"C0BFBDBB", x"BCBBB6B1", x"B2B3B1AC", x"A9A9A9A6",
									 -- x"A5A09F9F", x"9B999895", x"94908C88", x"87858280", x"7E7D7B77", x"726F6D6D", x"6C6A6663", x"6364625E",
									 -- x"5B5D5E5E", x"5C5A5857", x"54555655", x"524F4E4E", x"504C4849", x"4E504E4B", x"4B4D4F50", x"50515252",
									 -- x"52515153", x"5455585C", x"61605D5E", x"64656362", x"6566686A", x"6B6D7072", x"74737272", x"73757778",
									 -- x"787C7F80", x"7F7F8183", x"82848585", x"85878685", x"88898682", x"858B8880", x"82838587", x"87878888",
									 -- x"86858586", x"8787898A", x"888A8785", x"87858488", x"86858482", x"82848482", x"82848584", x"81808183",
									 -- x"807F7E80", x"82827F7C", x"7D79797A", x"78797A77", x"75757879", x"77747273", x"77726F6F", x"6F6D6A67",
									 -- x"706C696A", x"6C6D6A66", x"6969696A", x"6B696663", x"6A68645F", x"5E5F5F5E", x"5B5D5E5E", x"5C595857",
									 -- x"59575555", x"54525050", x"5050504E", x"4C4B4A4A", x"4D474242", x"4444413E", x"4443403F", x"3F3F3E3C",
									 -- x"BABAB9B8", x"B7B7B7B7", x"B6B7B8B8", x"B9BBBBB9", x"B6B7B8B8", x"B7B6B6B6", x"B1AFAEAE", x"ACA9A8A8",
									 -- x"A6A5A3A1", x"A1A3A2A0", x"A1A1A2A3", x"A19E9E9F", x"9E9C9D9E", x"9F9E9EA0", x"A4A5A7A9", x"ABABABAB",
									 -- x"AEADAAA6", x"A3A29D99", x"98979798", x"96939496", x"96979798", x"9B9E9F9E", x"A09E9C99", x"97989C9F",
									 -- x"A4A5A6A8", x"AEB3B4B2", x"B5B7B8B8", x"B8B9BABB", x"BFC0C1C2", x"C3C3C2C2", x"C3C2C4C7", x"CCCECECC",
									 -- x"C8C4C0BF", x"BEBDBEC0", x"C0C1C1C0", x"C0C0BDB9", x"B9B9B8B8", x"B8B9B9BA", x"BCBEC1C4", x"C4C4C6CA",
									 -- x"CBCCCCC9", x"CACDCCC8", x"C3C0BCBB", x"B9B7B5B6", x"B8B9B9B8", x"B8BBBCBB", x"B9BABBBB", x"BDBFBEBB",
									 -- x"BEBDBDBE", x"C0C2C4C5", x"C5C6C7C8", x"C8C6C4C3", x"C6C9CCCE", x"D0D0CECA", x"C5C5C4C3", x"C3C2C2C2",
									 -- x"C0BEBDBE", x"BFBEBFC0", x"C0C1C2C3", x"C2C3C4C5", x"C3C7CACA", x"CBCDCDCD", x"D0D1D2D3", x"D3D3D4D4",
									 -- x"D5D5D2CF", x"CECDCAC7", x"C8C6C4C4", x"C4C4C2C1", x"C2C3C4C4", x"C4C3C2C1", x"C1BFBEBE", x"C0C2C4C4",
									 -- x"C3C4C6C6", x"C6C5C4C3", x"C2C4C5C4", x"C2C3C4C4", x"C2C2C3C5", x"C7C7C9CC", x"CACBCED0", x"D3D4D4D3",
									 -- x"D4D4D5D5", x"D5D5D5D5", x"D7D8D9D9", x"DBDCDCDA", x"D8D9DDDC", x"D9DCDFDC", x"DDDDDCDC", x"DDDDDDDC",
									 -- x"DADAD9D7", x"D7D7D4D1", x"D2CFCAC5", x"C2C0C0C1", x"BFBDBBBA", x"B8B5B4B4", x"B2B3B0AB", x"A8A9A8A4",
									 -- x"A5A2A2A0", x"9C9C9A95", x"95918C89", x"88868481", x"81807E7A", x"7672706F", x"6A6A6866", x"65656361",
									 -- x"5E5F5F5D", x"5B5A5A5A", x"57575756", x"54514F4D", x"4F4C4A4C", x"50514D49", x"4B4B4C4D", x"4E505253",
									 -- x"50505154", x"56585B5E", x"5E5E5E5E", x"5F646764", x"6567696A", x"6B6D7072", x"75747272", x"73757778",
									 -- x"78797C7F", x"7E7C8086", x"82838482", x"82848484", x"84838281", x"83868581", x"82828283", x"84848483",
									 -- x"84838486", x"85838589", x"888A8481", x"85848083", x"82817F7D", x"7D80807F", x"81818181", x"81807E7D",
									 -- x"7D7C7B7B", x"7C7C7B7A", x"78757677", x"76777774", x"73727273", x"726F6C6C", x"716E6D6D", x"6C696868",
									 -- x"6A686667", x"69696764", x"67676869", x"69686564", x"67666461", x"6162615F", x"5D5E5E5C", x"5A585757",
									 -- x"59545152", x"53525050", x"4E4F4F4E", x"4C4A4948", x"45434141", x"4445423D", x"41403F3E", x"3D3D3D3D",
									 -- x"B8B8B7B7", x"B6B6B7B8", x"B9BABBBB", x"BCBDBDBB", x"B7B9BCBD", x"BBB9B8B8", x"B6B4B3B3", x"B1AEACAD",
									 -- x"ABACAAA7", x"A7AAA9A6", x"A6A4A3A2", x"9F9D9EA1", x"9B9A9B9E", x"9F9EA0A4", x"A7A6A6A9", x"ADAEADAC",
									 -- x"B0B0ADA8", x"A4A3A2A0", x"9A9A9A9A", x"97939395", x"9798999A", x"9DA0A09F", x"A0A09F9C", x"9A9B9EA1",
									 -- x"A4A5A6A8", x"ADB1B3B1", x"B5B6B9BB", x"BBBABABC", x"BDBEC0C1", x"C1C1C1C0", x"C0C1C3C5", x"C7C9CBCC",
									 -- x"CAC5C0BF", x"BEBDBFC2", x"C1C2C2C1", x"C1C1BEB9", x"BABAB9B8", x"B8B8B9BA", x"BDBEC1C4", x"C2C0C2C6",
									 -- x"C5C8C8C7", x"C8CBCAC5", x"C4C0BCBA", x"B8B5B4B3", x"B5B7B7B5", x"B5B7B8B6", x"B4B5B6B5", x"B7BBBCBB",
									 -- x"B8B7B6B7", x"BABCBDBD", x"C1C3C5C6", x"C5C4C4C4", x"C3C5C8CA", x"CCCCCAC7", x"C3C2C0BE", x"BDBDBEBE",
									 -- x"BDBDBDBD", x"BCBBBDC0", x"C0C1C2C2", x"C1C2C3C5", x"C1C5C9C9", x"CACCCDCD", x"D1D2D3D4", x"D4D4D5D6",
									 -- x"D5D6D4D0", x"CDCCCBCA", x"C9C7C5C4", x"C4C3C1C0", x"C2C3C4C4", x"C4C3C1C0", x"C1BFBCBB", x"BDBFC0C1",
									 -- x"C8C7C6C6", x"C6C4C1BE", x"C3C5C5C3", x"C2C4C2BF", x"C3C2C4C6", x"C7C6C8CB", x"CDCDCDCF", x"D1D3D5D5",
									 -- x"D4D3D3D4", x"D6D6D5D4", x"D4D7DADA", x"DADBDBD9", x"D9DBDFDD", x"D9DBDEDC", x"DFDEDDDD", x"DEDFDEDD",
									 -- x"D9DBDBD9", x"D8D7D4D1", x"CFCDCBC8", x"C5C4C3C3", x"BCBAB9B8", x"B4B0B1B6", x"B2B3B0AB", x"A9AAA8A4",
									 -- x"A5A4A4A2", x"9E9E9C94", x"94918C8A", x"89878482", x"7E7D7B79", x"76747271", x"6A6C6D6A", x"68686665",
									 -- x"62615F5C", x"59595A5C", x"59585655", x"54514D49", x"484A4C4E", x"4D4B4947", x"4E4D4B4A", x"4A4B4E50",
									 -- x"53535558", x"59595A5C", x"5D5D605E", x"5C656B66", x"67686B6C", x"6D6E7072", x"74727170", x"71747677",
									 -- x"7B797A7D", x"7A757981", x"7E7F7F7D", x"7C7E8080", x"807D7D7F", x"81807F81", x"80807F80", x"81818180",
									 -- x"82838586", x"84818387", x"8788807D", x"84837E7F", x"81807D7B", x"7C7E7F7E", x"7D7B7A7C", x"7E7E7975",
									 -- x"7B7A7877", x"76777777", x"74717273", x"7272736F", x"706D6C6F", x"706F6D6B", x"65666869", x"6765666A",
									 -- x"65656566", x"67666463", x"64646666", x"65646261", x"65666562", x"60605E5A", x"5D5D5D5B", x"5A585757",
									 -- x"59545050", x"51514F4D", x"4A4B4B4B", x"49474645", x"4343413F", x"4043413C", x"3D3D3D3C", x"3B3B3C3C",
									 -- x"BAB9B8B8", x"B9B9B9B8", x"B6B9BAB9", x"BABEC1C2", x"C0BFBFBF", x"BFBFBEBE", x"B9BBBCBA", x"B9B7B5B2",
									 -- x"B3B1AFAE", x"AEAFB0B0", x"ACA7A5A5", x"A39E9B9D", x"9C9B9B9E", x"A0A2A6A9", x"A4A8ACAE", x"AFB0B0AF",
									 -- x"AEADACAB", x"A9A6A3A0", x"9F9E9B98", x"95939290", x"92959697", x"9A9FA09E", x"A0A09E9D", x"9D9EA0A2",
									 -- x"A4A7A7A7", x"ABADAFB3", x"B2B6BBBC", x"BAB9BABB", x"BFBFBFBF", x"BFC0C1C2", x"C5C4C2C0", x"C3C9CBCA",
									 -- x"C9C7C4C2", x"C1C1C2C3", x"C2C3C3C2", x"C0BEBDBD", x"BFBBB7B6", x"B7B9B8B7", x"BBBBBEC1", x"C1C0BFC1",
									 -- x"C4C3C2C4", x"C6C8CBCD", x"C2BDB9B7", x"B6B3B1B0", x"B0B3B4B1", x"B0B1B1B0", x"B3B0AFB0", x"B3B4B3B1",
									 -- x"B1B2B1AE", x"B0B4B4B0", x"BABABBBD", x"BFC0C0C0", x"BFC3C4C2", x"C3C7C7C5", x"C4C1BFBE", x"BCBABBBD",
									 -- x"BABBBCBB", x"BBBBBCBD", x"BCBEC1C2", x"C1C0C1C2", x"C2C4C8CA", x"CBCCCCCC", x"D3D0D2D6", x"D8D5D4D5",
									 -- x"D4D3D1D0", x"CFCDCCCB", x"CCC8C5C4", x"C6C6C4C2", x"C2C2C3C5", x"C3C1C2C4", x"C1C2C1BF", x"BDBFC0C0",
									 -- x"C7C6C5C4", x"C4C3C2C1", x"C2C0C0C2", x"C2C1C2C4", x"C0C2C4C6", x"C7C6C6C6", x"C8CED0CD", x"CFD5D7D3",
									 -- x"D4D3D3D4", x"D3D1D2D5", x"D7D7D8DB", x"DCDADADA", x"DBDDDEDD", x"DDDFE0E0", x"E0DFDEDE", x"DEDEDEDE",
									 -- x"DBDBDBD9", x"D6D3D2D2", x"CDCBC9C7", x"C4C3C1C0", x"BEBABDB9", x"B3B0AFB6", x"B0AEABAA", x"A9A7A6A6",
									 -- x"A2A6A59E", x"9B9C9B97", x"8F8F8D8B", x"88848281", x"79797B79", x"73717270", x"706B696B", x"69646469",
									 -- x"615D5B5B", x"5B575554", x"5E575253", x"53504F51", x"4E4F4E4C", x"4F54524B", x"504D4B4B", x"4C4E5357",
									 -- x"53525255", x"56585B5E", x"5A636763", x"60636665", x"6467676A", x"6F717072", x"6D72736F", x"70757671",
									 -- x"7877787A", x"7A7A7C80", x"807F807F", x"7E7F807B", x"7F7D7C7D", x"7E7D7C7C", x"7B7E7F7D", x"7B7D7F7F",
									 -- x"81807F7F", x"7F7F7F7E", x"82828281", x"7E7C7C7F", x"807C7C7C", x"78787A79", x"79777575", x"77787776",
									 -- x"74737273", x"73717070", x"7372706E", x"6C6C6E6F", x"6E67666D", x"6E69696D", x"65696864", x"6467655F",
									 -- x"5E5F6161", x"61626364", x"60626569", x"69656261", x"60636664", x"615F6062", x"5E5B5A5B", x"5B585350",
									 -- x"534F4D4F", x"514F4C4B", x"4F4B4848", x"48454545", x"43403E3F", x"3E3D3D3E", x"3E3B3B3D", x"3C393535",
									 -- x"BAB9B8B8", x"B9BABBBB", x"B9BCBDBC", x"BCC0C3C4", x"C3C2C1C1", x"C1C2C3C3", x"C2C3C3C1", x"C0BFBEBC",
									 -- x"B5B3B2B4", x"B5B5B1AE", x"ADABA7A3", x"A09F9E9D", x"9E9C9D9F", x"A1A3A6A9", x"AAADAFB0", x"B0B0AFAD",
									 -- x"B0AFAEAC", x"AAA6A29F", x"9F9E9C99", x"96949292", x"91939596", x"999D9F9E", x"9F9F9F9F", x"9FA0A2A3",
									 -- x"A4A7A6A6", x"AAACAEB2", x"B1B4B8B9", x"B9B9BBBC", x"BCBDBEBF", x"C0C0C1C1", x"C0C2C3C2", x"C3C7C9C9",
									 -- x"CBC7C3C1", x"C2C4C4C4", x"C5C5C5C4", x"C2C0BFBF", x"BEBCBAB9", x"BABAB9B7", x"B7B8BBBE", x"BFBEBEBF",
									 -- x"BFC0C3C6", x"C8C8C8C7", x"C5BFBAB7", x"B5B1AEAD", x"ADAFAFAE", x"ADADADAC", x"AFADACAE", x"B0B1AFAD",
									 -- x"B0AFADAA", x"AAACAFAF", x"B2B2B3B4", x"B4B7BABD", x"C0BEBEBF", x"C1C2C3C3", x"C1BEBBBA", x"B9B7B6B6",
									 -- x"B6B8B9B9", x"B8B8B9BA", x"BDBDBEBF", x"C0C1C1C1", x"C4C4C5C6", x"C6C8CACB", x"CDCFD1D2", x"D4D5D5D5",
									 -- x"D3D2D1D0", x"D0CFCDCC", x"CCCAC7C6", x"C6C5C4C3", x"C3C3C3C4", x"C3C0C0C1", x"C0C1C1BF", x"BEC0C1C1",
									 -- x"C2C2C2C2", x"C2C1BFBE", x"C2C0BFC0", x"C0BEBEC0", x"C1C3C5C6", x"C7C7C8C8", x"C7CCCFCF", x"D0D3D3D1",
									 -- x"D2D2D3D5", x"D4D3D4D7", x"D6D5D6D8", x"D9D8D9DA", x"DADCDCDB", x"DBDDDEDE", x"E0DFDEDE", x"DEDFDEDE",
									 -- x"DADADAD9", x"D7D5D4D3", x"CECECDCA", x"C5C1BFBE", x"BEBBBCB8", x"B5B4B1B5", x"B2AFACAC", x"ACAAA8A7",
									 -- x"A7A5A29F", x"9D9B9895", x"92918F8B", x"88858382", x"7E7C7D7B", x"75737371", x"6D6C6A68", x"66646465",
									 -- x"62605F5F", x"5D595757", x"5D575354", x"54514F4F", x"4D4C4C4D", x"4E4E4F52", x"4F4D4C4D", x"4E4E5053",
									 -- x"51525456", x"5555585C", x"5A5F605C", x"5C626766", x"6A6B6766", x"6A6D7075", x"72737370", x"71757674",
									 -- x"7575787A", x"7B7A7C7F", x"807F7F7D", x"787A7D7C", x"797B7C7B", x"7978797A", x"787B7D7C", x"7B7C7C7C",
									 -- x"7E7E7D7D", x"7D7C7C7C", x"7C7F7F7B", x"78797A79", x"7877797A", x"76767672", x"78767474", x"74747270",
									 -- x"75737070", x"6E6C6B6B", x"6D6C6B69", x"68696B6C", x"66646469", x"6B696665", x"68696763", x"6263625E",
									 -- x"61616261", x"60606061", x"5D636766", x"65656563", x"62646462", x"5F5D5E5F", x"5C5B5959", x"59595755",
									 -- x"57524F4F", x"4F4D4B4B", x"4B484647", x"47454444", x"42403F40", x"3F3E3D3D", x"3D3B3C3E", x"3D393534",
									 -- x"BCBBB9B9", x"B9BABBBB", x"BCBEBFBE", x"BFC1C4C5", x"C6C5C4C3", x"C4C6C8C9", x"C9C9C8C5", x"C4C4C4C2",
									 -- x"BAB8B7B9", x"BBBAB5B0", x"B0B0ABA2", x"A0A2A29E", x"9C9B9CA0", x"A3A6A9AC", x"B0B1B2B1", x"B1B1AFAC",
									 -- x"B0AFAFAD", x"AAA6A19E", x"9D9D9C9A", x"97949394", x"91939495", x"989C9FA0", x"9E9FA0A1", x"A2A2A2A2",
									 -- x"A3A6A5A5", x"A9ABADB1", x"B2B4B6B7", x"B8BABCBD", x"BABBBDC0", x"C1C1C0BF", x"BEC1C4C4", x"C4C6C9CA",
									 -- x"CBC6C1C0", x"C3C6C6C5", x"C7C7C7C6", x"C4C2C1C0", x"BDBDBDBC", x"BBB9B8B7", x"B7B8BABE", x"BFBDBEBF",
									 -- x"BBBDC1C4", x"C5C5C4C3", x"C5BFB9B6", x"B3AFACAA", x"ACACACAB", x"ABACABA9", x"AAA8A8A9", x"ABABA9A7",
									 -- x"ADACACAA", x"A8A7AAAD", x"ABADAFAF", x"AEB0B4B8", x"BDB7B4B9", x"BCBCBCBF", x"BCB9B7B7", x"B8B6B3B2",
									 -- x"B4B6B7B7", x"B7B6B7B8", x"BDBBBABB", x"BEC0C0BF", x"C3C3C3C3", x"C3C4C6C7", x"C7CDD0CF", x"D0D4D4D2",
									 -- x"D0D0CFCF", x"D0CFCECD", x"CAC9C8C7", x"C5C4C4C4", x"C5C3C3C4", x"C4C2C0C0", x"C2C4C3C1", x"C0C2C3C3",
									 -- x"C0C1C2C3", x"C3C1BFBE", x"C0BFBFC0", x"BFBEBDBE", x"C1C3C4C6", x"C7C8C9CA", x"C9CACDCE", x"CFCFD0D0",
									 -- x"D1D2D4D5", x"D5D4D5D7", x"D5D4D3D4", x"D5D5D7DA", x"D9DBDCDB", x"DBDDDEDE", x"DFDEDEDF", x"DFDFDEDE",
									 -- x"DCDBD9D9", x"D8D7D5D3", x"CECFD0CD", x"C6C1BEBE", x"BEBBBCB6", x"B4B6B1B1", x"B1ADAAAB", x"ACAAA7A6",
									 -- x"AAA4A0A1", x"A19D9896", x"9694908C", x"88858483", x"837F7F7D", x"77767572", x"6E6F6E69", x"67676663",
									 -- x"61616161", x"5E5B5A5C", x"5D585658", x"58545151", x"514C4D50", x"4D484B55", x"4E4C4B4E", x"4F4F4E4F",
									 -- x"51535556", x"5454585D", x"5C5E5D59", x"5A626969", x"6A6E6E6D", x"6E6E6E73", x"74727070", x"71737577",
									 -- x"7374777A", x"7B7A7B7C", x"7C7D7F7C", x"75757A7A", x"777A7A78", x"77787977", x"76797A7B", x"7B7C7A78",
									 -- x"797A7B7A", x"7978797A", x"787D7D77", x"74787874", x"72737675", x"7274736E", x"74727170", x"706E6B69",
									 -- x"6F6C6A6A", x"6A69696A", x"69686766", x"66676869", x"67656260", x"63666663", x"67666462", x"6161605F",
									 -- x"5E5F5F5F", x"60606162", x"5F676B66", x"63666765", x"65636260", x"5E5D5D5D", x"59595653", x"53565755",
									 -- x"5754504F", x"4F4D4B4B", x"4A484747", x"47464545", x"413F3F40", x"403E3C3C", x"3A3A3A3B", x"3A383839",
									 -- x"BEBDBBBA", x"BABABAB9", x"BDBFC1C0", x"C0C3C6C7", x"C7C7C6C6", x"C7C9CCCE", x"CCCCCBC7", x"C5C5C4C2",
									 -- x"C0BEBBBB", x"BCBCBAB7", x"B6B4AEA7", x"A3A3A2A0", x"9D9C9DA0", x"A3A5A8AB", x"B0B1B1B0", x"B1B2B0AE",
									 -- x"ADADADAC", x"AAA5A09D", x"9A9A9A99", x"96939395", x"92939496", x"989CA0A2", x"A0A0A1A2", x"A2A2A1A0",
									 -- x"A3A5A4A4", x"A8AAABB0", x"B3B3B3B4", x"B6B8B9BA", x"BABBBDBF", x"C0C0C0BF", x"BFC1C3C5", x"C6C8C9CB",
									 -- x"C9C6C2C0", x"C2C6C7C7", x"C8C8C8C7", x"C4C2C1C1", x"BCBDBDBC", x"BAB8B7B7", x"B8B8BBBE", x"BEBDBDBE",
									 -- x"B9BBBDBE", x"BFC1C2C2", x"C1BCB6B3", x"B1AEABAA", x"ABAAA9A8", x"A9A9A7A5", x"A5A4A3A3", x"A5A6A5A4",
									 -- x"A9A8A9AC", x"AAA7A6A9", x"A8AAADAE", x"AEAEAFB0", x"B3B0AFB2", x"B4B4B5B7", x"B5B2B0B2", x"B5B4B2B1",
									 -- x"B2B4B5B6", x"B5B5B6B7", x"BBB9B8B8", x"BABDBEBF", x"C0C2C3C3", x"C3C3C3C3", x"C5CBCFCF", x"CECFCFCD",
									 -- x"CDCDCDCE", x"CECECCCB", x"C7C7C6C6", x"C5C5C5C5", x"C5C4C4C5", x"C6C5C3C2", x"C4C5C4C2", x"C1C2C2C2",
									 -- x"C1C2C3C3", x"C2C0BFBE", x"BFBFBFC1", x"C1C0C0C0", x"C1C2C4C6", x"C7C8C9CA", x"CBC9C9CB", x"CCCBCED2",
									 -- x"D0D2D4D5", x"D5D4D4D5", x"D5D3D2D3", x"D4D4D6D9", x"DADCDDDD", x"DDDEDFDF", x"DEDEDEDF", x"DFDFDEDD",
									 -- x"DEDCDAD9", x"D9D8D4D1", x"CECECECC", x"C7C3C0BF", x"BCBBBCB5", x"B2B5AFAE", x"B1ACA8A8", x"AAA9A7A5",
									 -- x"A5A29FA0", x"A19F9A97", x"9895908B", x"88868685", x"847F7E7D", x"78777774", x"70706F6C", x"6A686664",
									 -- x"6261605F", x"5E5E5E5E", x"5B585758", x"59565454", x"534E4D50", x"4F4B4D54", x"504D4C4E", x"51515050",
									 -- x"53535453", x"5253595F", x"5B5E5E5A", x"5B626769", x"686E7171", x"706D6C70", x"726E6C6E", x"70717376",
									 -- x"73757879", x"79787879", x"777A7E7C", x"76757775", x"78787674", x"777A7872", x"74757677", x"78787775",
									 -- x"75777978", x"76757778", x"77797975", x"73757573", x"7170716E", x"6B70726E", x"6D6C6C6B", x"6B6A6867",
									 -- x"69676667", x"68686869", x"68676564", x"64656666", x"66635F5E", x"61636361", x"61606061", x"62626364",
									 -- x"60616162", x"63646666", x"666A6A67", x"64656666", x"66636060", x"615F5E5E", x"59595550", x"51555551",
									 -- x"53525151", x"4F4D4B4A", x"49484646", x"45444343", x"403F3E3F", x"3F3C3A3A", x"3B3A3937", x"3535383A",
									 -- x"BEBDBCBC", x"BBBBBAB9", x"BEC0C2C2", x"C3C6C8C9", x"C9C9CACB", x"CBCDCFD0", x"D1D1D0CC", x"C9C8C6C3",
									 -- x"C2C1BFBE", x"BDBCBDBD", x"BBB6B1AD", x"A9A3A0A0", x"A09F9E9F", x"A0A1A3A5", x"ADAEAFAE", x"AFB1B0AE",
									 -- x"ADADADAD", x"AAA5A09C", x"97969697", x"95929395", x"92939496", x"989B9FA2", x"A0A0A0A1", x"A2A2A2A1",
									 -- x"A3A5A5A5", x"A9AAABAF", x"B1B1B1B1", x"B3B5B7B8", x"BBBCBDBF", x"C0C0C0C0", x"C1C0C1C3", x"C6C8CACA",
									 -- x"C7C8C5C2", x"C1C5C9CA", x"C9C9C9C7", x"C5C3C2C1", x"BDBEBDBB", x"B8B7B7B8", x"B8B8BABC", x"BCBAB9BA",
									 -- x"B8BBBCBB", x"BCBFC1C0", x"BEB9B4B2", x"B1AEABAB", x"A8A6A5A5", x"A5A4A2A1", x"A3A2A0A0", x"A1A3A3A3",
									 -- x"A6A3A4A8", x"A9A6A5A6", x"A7A7A8AA", x"ABACABA9", x"ABAFB0AE", x"AEAFB0AF", x"AFABA9AB", x"AFAFAEAE",
									 -- x"AEB0B1B2", x"B1B1B3B4", x"B7B8B8B8", x"B8BBBEC1", x"C0C1C2C2", x"C1C1C2C2", x"C4C6CBCF", x"CECAC9CB",
									 -- x"CDCCCCCC", x"CDCCCBCA", x"C8C7C5C6", x"C7C7C6C5", x"C5C5C4C5", x"C6C6C4C2", x"C3C4C3C1", x"C0C0C1C0",
									 -- x"C2C2C2C1", x"BFBEBEBF", x"BEBFC0C1", x"C1C2C2C2", x"C2C4C6C8", x"C9C9C9CA", x"CAC7C7CA", x"CACACDD2",
									 -- x"CDD0D3D4", x"D4D4D5D5", x"D5D3D3D4", x"D5D5D6D8", x"DADCDDDD", x"DDDFDFDF", x"DEDEDEDE", x"DFDFDEDD",
									 -- x"DEDCD9D9", x"D9D8D4D1", x"CFCDCAC8", x"C6C4C1BE", x"BCBCBEB6", x"B1B2AEAD", x"B1ACA7A7", x"A9A9A7A6",
									 -- x"9EA1A19D", x"9D9E9B96", x"97948F8B", x"88878787", x"817D7D7C", x"78787975", x"706C6B6E", x"6D696768",
									 -- x"67645F5E", x"5F61605F", x"57555455", x"56565656", x"524E4B4D", x"50525150", x"534F4C4E", x"50525354",
									 -- x"53525253", x"5353565A", x"575D605E", x"5C5E6264", x"676C6D6B", x"6A696A70", x"6F6A696D", x"6F6F7073",
									 -- x"72747676", x"75757677", x"75767A7A", x"76777773", x"74757472", x"72757470", x"71717172", x"72727271",
									 -- x"72747676", x"74747576", x"76737374", x"726F6F72", x"6F6E6D6A", x"676C6F6C", x"6A696867", x"67676767",
									 -- x"69676666", x"66646263", x"65636161", x"61626262", x"5F5D5F64", x"65605B5A", x"5C5C5F63", x"66666769",
									 -- x"6B6B6B6B", x"6B6B6B6B", x"6D696768", x"67656567", x"66626061", x"62605D5C", x"5C5A5552", x"54575550",
									 -- x"5151514F", x"4D4C4B4A", x"47474442", x"403F3F3F", x"403E3D3D", x"3C3A3939", x"3C3C3A36", x"33323334",
									 -- x"BEBDBCBC", x"BCBDBCBC", x"BFC2C4C4", x"C5C8CBCB", x"CBCDCFCF", x"CFD0D1D2", x"D2D3D2CF", x"CDCBC8C5",
									 -- x"C3C4C4C3", x"C1BFBEBF", x"BEB8B4B2", x"ADA5A0A1", x"A09E9D9E", x"A0A1A4A7", x"ABADAEAD", x"ADAEAEAE",
									 -- x"AFAFAFAE", x"ABA5A09C", x"97949395", x"94929294", x"92929395", x"96989CA1", x"9F9E9EA0", x"A2A4A4A4",
									 -- x"A3A6A6A7", x"AAABABAF", x"B0B0B2B3", x"B4B6B8BA", x"BCBCBDBE", x"BFBFC0C0", x"C2BFBFC2", x"C5C7C8C9",
									 -- x"C8CAC8C4", x"C2C6CACB", x"CACACAC8", x"C6C4C2C2", x"BEBEBDBA", x"B8B7B8BA", x"B8B8BABB", x"BAB7B6B7",
									 -- x"B5B9BCBA", x"BABCBCBB", x"BBB7B3B1", x"B0AEABAA", x"A6A5A4A4", x"A3A1A0A0", x"A1A09F9F", x"A0A2A3A3",
									 -- x"A6A3A1A3", x"A5A6A7A7", x"A8A5A4A5", x"A8AAAAA8", x"A8AFB1AE", x"ABACACA9", x"ACA9A7A8", x"AAABAAAA",
									 -- x"ACADAEAE", x"AEAFB1B2", x"B4B5B7B7", x"B8BABEC1", x"C2C1BFBE", x"BEBFC2C4", x"C2C2C6CC", x"CCC8C6C9",
									 -- x"CDCCCBCB", x"CBCBCACA", x"CAC9C7C7", x"C8C7C6C4", x"C5C5C4C3", x"C3C4C3C1", x"C3C4C4C2", x"C1C2C3C2",
									 -- x"C3C3C2C0", x"BEBDBFC0", x"BEBFC0BF", x"C0C1C1C0", x"C5C6C8C9", x"C9CACACA", x"C7C6C8CB", x"CCCACBCE",
									 -- x"CACED2D3", x"D4D6D7D7", x"D7D5D5D6", x"D6D6D6D8", x"D8DADCDC", x"DCDEDEDD", x"DEDEDDDD", x"DEDEDDDC",
									 -- x"DCDAD8D8", x"D9D8D5D2", x"D1CDC9C6", x"C5C4C0BD", x"BEBDBFB7", x"B2B2AEB0", x"AFAAA6A6", x"A7A6A5A4",
									 -- x"9EA4A5A0", x"9D9E9C96", x"96938E8B", x"8A898887", x"7F7D7D7C", x"79787977", x"716C6B71", x"726D6B6E",
									 -- x"6E69635F", x"6163625E", x"57565656", x"57585858", x"54534E4B", x"4F545047", x"504C494A", x"4C4E5154",
									 -- x"54535456", x"56545455", x"575D6261", x"5E5E6062", x"62686B6B", x"6B69686D", x"6C69686B", x"6E6E6F70",
									 -- x"6F717271", x"71737575", x"75737474", x"73767672", x"6F727573", x"6F6D7073", x"72717070", x"706F7071",
									 -- x"6F717373", x"72727373", x"75706F72", x"716C6C70", x"6E6B6D6D", x"6A6A6B69", x"69686765", x"65646565",
									 -- x"66646364", x"63615F5F", x"61605E5E", x"60616161", x"5E5C5F64", x"645E5B5D", x"5C5F6468", x"6A6B6C6C",
									 -- x"6F6F6F70", x"71717170", x"716A686B", x"6C68676B", x"66615F61", x"625E5B5A", x"5B585454", x"55565451",
									 -- x"5353514D", x"4A494A4B", x"46464541", x"3F3F3F3F", x"403E3C3C", x"3C393839", x"37383836", x"35333230",
									 -- x"C0BFBDBC", x"BDBEBFBF", x"C0C3C5C5", x"C6C8CBCB", x"CDCED0D1", x"D0D0D1D3", x"D1D2D1CF", x"CDCCCAC7",
									 -- x"C7C7C7C6", x"C5C3C0BF", x"C0BDB9B6", x"B1AAA5A3", x"A09E9D9E", x"A0A2A6AA", x"A9ADAFAE", x"ACACADAD",
									 -- x"AFAFAEAD", x"AAA5A09D", x"9B959294", x"94929193", x"92929396", x"96979BA0", x"9F9E9EA1", x"A4A6A6A5",
									 -- x"A4A8A8A9", x"ADADACAF", x"AFB1B4B5", x"B5B6B8BA", x"BBBBBCBD", x"BEBFC0C0", x"C1C0C0C3", x"C5C6C7C9",
									 -- x"C8CAC8C3", x"C2C6C9C8", x"CACACAC8", x"C5C3C1C1", x"BDBCBBB9", x"B8B7B8B8", x"B7B7B8BA", x"B8B5B4B4",
									 -- x"B2B7B9B6", x"B5B6B6B4", x"B5B1AFAF", x"AEACA9A8", x"A5A4A4A4", x"A29F9EA0", x"9C9C9D9E", x"9F9FA0A0",
									 -- x"A3A3A2A1", x"A2A5A7A7", x"A6A5A4A4", x"A6A7A6A6", x"A7A9ACAC", x"ABAAA9A9", x"A9A7A6A8", x"A8A7A6A7",
									 -- x"A9AAABAA", x"AAABAEB0", x"B0B1B2B4", x"B7BABCBE", x"C1C0BEBC", x"BBBDC0C2", x"BFC0C3C6", x"C7C7C7C7",
									 -- x"CBCAC8C8", x"C8C9C9C9", x"C8C8C8C7", x"C6C5C4C4", x"C3C5C5C3", x"C2C3C4C3", x"C3C5C5C3", x"C2C3C3C2",
									 -- x"C2C2C1BF", x"BDBDBFC1", x"BEC0C0BF", x"BFC1C2C0", x"C8C8C8C7", x"C7C8C9CA", x"C7C8C9CB", x"CBCBCBCC",
									 -- x"CACED2D2", x"D4D6D8D8", x"D9D7D7D7", x"D7D6D7D8", x"D6D9DBDB", x"DBDDDDDC", x"DFDEDDDC", x"DCDCDCDB",
									 -- x"DAD9D7D7", x"D8D7D4D2", x"D0CECAC7", x"C5C3C0BE", x"C1BBBCB7", x"B4B3AFB1", x"ACA9A6A6", x"A5A3A2A2",
									 -- x"A0A4A5A3", x"9F9D9B98", x"96938F8C", x"8B8A8987", x"817F807F", x"7A797A78", x"75717072", x"73716F6F",
									 -- x"6E6B6763", x"63646360", x"5B5B5A5A", x"5A5A5A59", x"5757534E", x"4E504D47", x"4C4A494A", x"4B4C4F53",
									 -- x"51525354", x"53525456", x"595D605F", x"5E5F6264", x"5E65696B", x"6D6A676A", x"6B696769", x"6B6D6D6C",
									 -- x"6B6E6F6E", x"6E6F7171", x"716F7171", x"7073736F", x"6F6E7071", x"6E6B6C71", x"72717070", x"6F6D6E70",
									 -- x"6C6D6E6F", x"7070706F", x"716E6D6E", x"6D6B6A6C", x"6C68696D", x"69656564", x"65656462", x"61605F5F",
									 -- x"5F5D5D5E", x"5F5E5D5E", x"5F5D5B5C", x"5D5E5E5D", x"5F5F5E5E", x"5C5D6064", x"61676B6C", x"6E70716F",
									 -- x"6D6E6F71", x"73747372", x"716E6C6D", x"6D6A696B", x"66615F61", x"625E5B5C", x"59565455", x"54515153",
									 -- x"5254534F", x"4A494949", x"43454643", x"41414140", x"403E3D3E", x"3D3A3838", x"35363634", x"34353431",
									 -- x"C4C2BEBC", x"BCBEC0C1", x"C0C3C5C5", x"C5C7C9C9", x"CDCFD0D0", x"CFCFD0D2", x"D0D1D1CF", x"CECECDCB",
									 -- x"CCCAC8C6", x"C6C5C3C0", x"C2C2BFB8", x"B3B0ABA5", x"A6A3A0A0", x"A0A1A4A7", x"A7ACB0AF", x"ACACAEAF",
									 -- x"ADACACAB", x"A9A5A19D", x"9E979394", x"95939293", x"93939597", x"98989BA0", x"A09FA0A2", x"A5A7A6A4",
									 -- x"A4A8A9AB", x"AEAEADAF", x"ADB0B4B4", x"B3B2B4B6", x"B8B9BBBD", x"BEBFBFC0", x"C1C1C3C6", x"C6C5C7CA",
									 -- x"C8C9C6C1", x"C2C6C7C4", x"C8C9C8C6", x"C4C1C0BF", x"BBBAB9B8", x"B7B7B6B6", x"B3B3B5B6", x"B4B1B0B0",
									 -- x"B1B5B5B0", x"AEAFB0AF", x"AFACAAAB", x"ACAAA7A6", x"A3A2A2A2", x"9F9C9B9D", x"97989A9C", x"9D9D9C9C",
									 -- x"9CA0A2A0", x"A0A2A4A2", x"A2A3A4A5", x"A4A2A1A0", x"A5A3A5AA", x"ACA9A9AB", x"A3A3A4A6", x"A5A3A2A3",
									 -- x"A5A6A6A6", x"A6A7AAAC", x"ACACADB1", x"B5B9BABA", x"BEBEBDBC", x"BCBCBDBE", x"BFC1C2C0", x"C2C6C7C4",
									 -- x"C8C6C5C4", x"C5C6C7C7", x"C4C5C7C6", x"C4C2C3C4", x"C2C5C5C3", x"C2C4C6C6", x"C1C3C3C0", x"BFBFBFBE",
									 -- x"BEBEBEBD", x"BBBBBDBF", x"BFC0C0BF", x"C0C2C3C2", x"C9C8C6C4", x"C4C5C7C9", x"C9CACAC8", x"C8CACCCC",
									 -- x"CCD0D3D3", x"D4D6D8D8", x"DBD9D7D7", x"D7D6D7D9", x"D6D9DBDB", x"DBDDDDDC", x"DFDEDCDC", x"DBDBDBDB",
									 -- x"DBD9D8D7", x"D6D5D2D0", x"CECDCBC8", x"C5C2C1C0", x"C1B9B8B6", x"B5B4AEB1", x"ACAAA9A9", x"A8A4A2A2",
									 -- x"A09FA0A2", x"9F9A9797", x"9693908D", x"8C8B8987", x"83828482", x"7C797A78", x"77767471", x"70706E6A",
									 -- x"6B6B6865", x"64656461", x"5D5D5D5B", x"5B5A5957", x"55555451", x"4F50504F", x"4D4D4D4E", x"4F4F5154",
									 -- x"4D4D4E4D", x"4B4C5259", x"5A5B5B5A", x"5B5E6264", x"61656463", x"6566676C", x"6B696666", x"686B6B69",
									 -- x"6A6D6E6C", x"6B6C6D6C", x"6B6C7072", x"7071706A", x"7068666B", x"6E6B6869", x"6E6E6E6E", x"6C68696D",
									 -- x"6A6A6B6D", x"6E6E6E6D", x"6B6B6A68", x"67686866", x"69626367", x"635E5E60", x"60606160", x"5E5C5B5A",
									 -- x"5D5B595A", x"5B5A5A5C", x"5C5A5858", x"59595856", x"565C5F5B", x"595D6060", x"656C706F", x"70747471",
									 -- x"71717274", x"75757371", x"6D6F6E6B", x"68676766", x"67625F62", x"625F5E60", x"5A575759", x"554E5056",
									 -- x"4E535553", x"4E4C4946", x"3F424443", x"4242413F", x"3F3E3E3F", x"3E3B3837", x"3D3B3631", x"31323230",
									 -- x"C7C4C1C0", x"C0C1C0C0", x"C1C2C4C5", x"C6C7C9CB", x"CECDCED0", x"D1CFD0D2", x"D1D0D0D0", x"D0CFCDCB",
									 -- x"CBCBCAC8", x"C5C3C2C3", x"C2C5C4BD", x"B6B2ADA8", x"A3A2A0A0", x"A1A2A2A2", x"A6AAADAD", x"ACADAEAE",
									 -- x"B0ADABAA", x"ABAAA5A1", x"A19B9593", x"93929292", x"9695979A", x"9B9A9C9F", x"9CA0A4A5", x"A4A4A6A9",
									 -- x"A9AAABAB", x"ABADAEB0", x"ADB0B2B3", x"B3B4B6B9", x"BABBBDBE", x"BEBEBEBF", x"C3C2C2C1", x"C2C4C6C8",
									 -- x"C6C7C6C3", x"C0C0C4C7", x"C7C8C7C5", x"C5C4C0BC", x"BAB9B8B7", x"B7B6B5B4", x"B7B6B4B3", x"B2B0AFAE",
									 -- x"AFB0B1B0", x"AFACABAA", x"ABAAA8A8", x"A7A5A4A2", x"A09D9E9D", x"98989A99", x"999A9997", x"97999A99",
									 -- x"9B9D9F9E", x"9FA2A4A4", x"A0A2A3A3", x"A2A1A1A1", x"A4A4A4A6", x"A8AAAAAA", x"A4A6A7A6", x"A4A3A3A5",
									 -- x"A4A4A4A4", x"A4A4A5A6", x"A7ADAFAC", x"AEB5B8B6", x"BDBCBAB9", x"BCBFBDB8", x"BEBEBDBE", x"BFC1C3C4",
									 -- x"C4C5C6C6", x"C4C3C4C5", x"C4C7C8C5", x"C3C4C4C3", x"C5C2C3C3", x"C0C2C5C3", x"C1C2C1BE", x"BFC2C1BC",
									 -- x"BBBBBBBC", x"BDBDBEBE", x"C1C0C0C2", x"C4C4C4C5", x"C7C5C4C6", x"C6C6C8CA", x"C8C8C8C7", x"CACCCCCA",
									 -- x"CED2D4D3", x"D4D9DBDA", x"D9DADBDA", x"D8D8D9DB", x"DADBDCDC", x"DCDBDCDC", x"DCDCDDDE", x"DEDDDCDC",
									 -- x"DBDAD8D7", x"D6D4D1CF", x"D1CECCCB", x"C7C1BFC0", x"BDB7B7B9", x"B5B0AEAD", x"AEAAA9AA", x"A8A3A2A4",
									 -- x"A29E9FA3", x"A19A999E", x"9493908D", x"8988898A", x"82878782", x"7E7D7D7B", x"7E767272", x"7375746E",
									 -- x"6E6C726A", x"676A6366", x"6262615F", x"5F5F5B56", x"57585754", x"53545351", x"55514E51", x"53525050",
									 -- x"4C4E5153", x"514F5155", x"5557595E", x"58636561", x"66626165", x"66636162", x"67656565", x"64676A68",
									 -- x"66696C6D", x"6C6C6D70", x"6D6B6A6C", x"6B676668", x"6B69696B", x"6B6A6B6E", x"676D716F", x"6B686663",
									 -- x"6B6A6866", x"67696B6C", x"6B6A6A6A", x"68646466", x"64646462", x"605F5F5F", x"5A5E605E", x"5A595959",
									 -- x"5556575A", x"5A575555", x"58585655", x"565A5E60", x"605B575A", x"60646666", x"66707479", x"70717178",
									 -- x"78777879", x"77747373", x"7172716D", x"6A696969", x"6667645F", x"5D5F5E5B", x"57575758", x"57555354",
									 -- x"53525050", x"4F4D4C4D", x"42454441", x"4042413E", x"3C3D3D3B", x"39373636", x"37333133", x"352F2C32",
									 -- x"CCC9C4C1", x"C0C0C0C0", x"C3C3C4C4", x"C4C5C7C9", x"CBCBCDCF", x"D0CFD0D3", x"D1D0CFCF", x"CFCFCDCC",
									 -- x"CCCCCCCA", x"C7C5C4C4", x"C3C5C5C0", x"B8B2AEAB", x"A6A5A3A2", x"A2A2A2A1", x"A1A5A8A9", x"AAABABAA",
									 -- x"AEACA9AA", x"ABAAA6A3", x"9F9A9593", x"93939393", x"95949698", x"98979799", x"9C9FA2A3", x"A3A4A7A9",
									 -- x"A9AAAAAB", x"ACADAFB0", x"AFB0B1B2", x"B3B4B6B8", x"BABBBCBD", x"BDBDBEBF", x"C0C0C1C1", x"C2C3C5C7",
									 -- x"C6C6C5C2", x"BFBFC1C4", x"C2C3C3C2", x"C1C0BCB9", x"B9B8B7B7", x"B6B6B4B3", x"B4B4B4B3", x"B2B0ADAA",
									 -- x"ACADAEAE", x"ADABA9A8", x"A8A7A6A5", x"A5A4A2A1", x"A19D9C9B", x"97989A99", x"99999795", x"96979694",
									 -- x"95999D9F", x"A0A09F9D", x"A2A1A1A2", x"A3A3A2A1", x"A2A2A2A3", x"A5A6A6A5", x"A4A5A6A5", x"A3A2A3A4",
									 -- x"A2A2A1A0", x"A0A1A3A5", x"A7A8AAAA", x"ACAEB1B1", x"B6B6B4B4", x"B6BABAB7", x"BCBBBBBB", x"BCBDC0C2",
									 -- x"C3C4C5C5", x"C5C5C5C5", x"C4C6C5C3", x"C1C2C2C1", x"C1BEC0C1", x"BFC2C5C3", x"C0C2C1BE", x"BEC0BEBA",
									 -- x"BDBDBDBC", x"BCBDBDBD", x"BFBEBEC1", x"C3C4C4C6", x"C6C6C7C7", x"C6C4C6C9", x"C9CACBCA", x"CACCCDCD",
									 -- x"CED1D5D7", x"D9DBDCDC", x"DBDCDCDB", x"DADADBDD", x"DADCDEDE", x"DCDBDCDE", x"DEDEDFDE", x"DEDCDBDA",
									 -- x"DBDAD8D6", x"D5D4D1CF", x"CDCBCAC9", x"C5C1BFC0", x"BDB6B6B7", x"B4B0AFAE", x"ADABAAA9", x"A8A5A3A3",
									 -- x"A4A2A1A1", x"A19F9D9C", x"9996938F", x"8C898785", x"86888782", x"80807F7D", x"7D787676", x"73747571",
									 -- x"7171736F", x"6B696362", x"66656360", x"5F5F5C57", x"58575452", x"53545250", x"4F4D4D4E", x"4F4E4E50",
									 -- x"514E4D4F", x"52525151", x"5357585D", x"5B63605C", x"63626365", x"66656565", x"64626363", x"62676B69",
									 -- x"64666868", x"68686A6C", x"6C6A6968", x"67666566", x"66656567", x"67656668", x"66696B69", x"68676562",
									 -- x"65656666", x"66656565", x"67656464", x"62616366", x"6363615E", x"5C5B5C5D", x"5C5B5958", x"595A5855",
									 -- x"53535456", x"57565758", x"55555555", x"56585A5B", x"5F5B5A5E", x"6367696B", x"75757478", x"797B7878",
									 -- x"7D7B7B7C", x"7B787574", x"72716F6E", x"6C696867", x"63656663", x"5F5D5B59", x"5B5A5A5B", x"5A565351",
									 -- x"53514F4F", x"4F4D4D4D", x"4A474443", x"43423F3D", x"3B3C3C3C", x"3B393735", x"38353031", x"34302D30",
									 -- x"D5D0CAC4", x"C1C0C1C1", x"C4C4C4C3", x"C3C3C5C6", x"C6C8CBCD", x"CDCDD0D3", x"D1D0CFCF", x"CFCFCFCE",
									 -- x"CECECECC", x"C9C6C5C4", x"C3C4C5C3", x"BCB4AFAF", x"ABA9A7A6", x"A5A4A2A0", x"A0A2A5A6", x"A8A9A8A6",
									 -- x"A9A7A5A5", x"A7A7A4A1", x"9D989494", x"94949393", x"96969799", x"99989899", x"9C9D9FA0", x"A2A4A6A8",
									 -- x"A7A8A9AA", x"ABADAEB0", x"AFAFAFB0", x"B1B3B5B6", x"BABBBCBC", x"BCBDBDBE", x"BEBFC0C1", x"C1C1C2C2",
									 -- x"C5C4C3C0", x"BEBDBEC0", x"BDBFC1BF", x"BEBDBBB8", x"B8B7B6B6", x"B5B5B3B2", x"B3B3B2B1", x"AFADABA9",
									 -- x"ABACAEAE", x"ACAAA9A8", x"A8A7A6A5", x"A4A4A3A2", x"A19D9B99", x"96989A99", x"96969494", x"96989793",
									 -- x"93979C9D", x"9E9E9D9A", x"A09E9D9F", x"A2A3A19F", x"9F9F9FA0", x"A1A2A1A0", x"A3A4A4A3", x"A1A1A2A3",
									 -- x"A09F9E9C", x"9C9EA1A4", x"A5A4A5A9", x"A9A8AAAD", x"AFAFAFAF", x"B1B5B6B6", x"B8B8B9B8", x"B8BABDBF",
									 -- x"C1C1C1C2", x"C3C3C2C1", x"C4C4C2C1", x"C1C2C2C0", x"C1BFC1C1", x"BFC0C3C1", x"C1C2C1BE", x"BEBFBEBA",
									 -- x"BFBFBEBD", x"BDBDBEBE", x"BEBDBDBF", x"C1C2C2C4", x"C4C5C8C8", x"C5C3C4C8", x"C8CBCDCB", x"CBCCCECF",
									 -- x"D0D1D4D8", x"DBDCDDE0", x"DDDEDEDE", x"DCDCDEDF", x"DADDE0DF", x"DCDBDDE0", x"E0DFDFDE", x"DCDBDADA",
									 -- x"DAD9D7D5", x"D4D3D0CE", x"CBCAC9C7", x"C4C0BEBE", x"BDB6B5B7", x"B3B0B0AE", x"AAABABA9", x"A7A6A4A2",
									 -- x"A6A6A3A0", x"A0A29F9A", x"97949290", x"908E8A87", x"88898681", x"8183827F", x"7D7B7C7B", x"76757775",
									 -- x"71747171", x"706C6C66", x"68676361", x"605F5D59", x"5B585351", x"53555451", x"4D4E5050", x"4E4D4F52",
									 -- x"534F4D4F", x"51525252", x"53585458", x"5A605958", x"5E606263", x"65676665", x"63616161", x"61656967",
									 -- x"64646363", x"63656668", x"68686663", x"62646464", x"61616364", x"64626263", x"65656463", x"64656361",
									 -- x"60626464", x"62616061", x"63616161", x"61606264", x"615F5C59", x"5757595A", x"5A585553", x"54565552",
									 -- x"54525152", x"52515254", x"52535455", x"55565859", x"5D5D6064", x"686B6F73", x"7A767576", x"7E81827E",
									 -- x"817E7D7F", x"7F7B7876", x"746F6D6E", x"6F6B6867", x"63656665", x"615B595A", x"5D5A595B", x"5C5A5756",
									 -- x"54504D4E", x"4E4D4C4C", x"4C454144", x"46424040", x"3C3B3B3C", x"3B393633", x"3836302F", x"32322E2D",
									 -- x"DAD6D0CA", x"C5C3C2C2", x"C4C4C4C3", x"C3C3C3C3", x"C3C5C8CA", x"CACBCDD0", x"D0D0D1D1", x"D1D1D1D0",
									 -- x"D0D0CFCD", x"CBC7C5C3", x"C3C3C4C4", x"BEB5B1B2", x"ADACAAA9", x"A8A7A4A1", x"A4A4A4A5", x"A7A8A6A4",
									 -- x"A5A3A1A2", x"A3A3A2A0", x"9C989594", x"94939292", x"96979899", x"9A9B9C9E", x"9D9D9D9E", x"A0A3A4A5",
									 -- x"A5A6A8A9", x"AAABADAF", x"AFAEADAE", x"AFB1B3B3", x"B9BABCBD", x"BDBCBDBD", x"BFBFC0C0", x"BFBFBFBF",
									 -- x"C2C2C0BE", x"BDBCBCBC", x"BBBEC0BF", x"BDBCBBBA", x"B6B5B5B4", x"B4B3B1B0", x"B4B1AEAC", x"ABABABAB",
									 -- x"AAABABAB", x"AAA9A8A8", x"A8A7A5A4", x"A3A2A2A1", x"A19C9A99", x"97989B98", x"96969695", x"96989795",
									 -- x"97999B9B", x"9B9D9E9D", x"9D9C9C9D", x"A0A1A19F", x"9D9E9E9F", x"9F9F9F9E", x"A1A2A3A2", x"A1A0A0A1",
									 -- x"9F9E9D9B", x"9B9C9FA1", x"A2A2A4A7", x"A8A7A8AB", x"ACADADAE", x"AFB2B4B5", x"B4B6B7B8", x"B8B9BBBE",
									 -- x"C0BFBFBF", x"C0C0BEBD", x"C3C2C1C1", x"C2C3C2C0", x"C0BEBFC0", x"BEBFC1BE", x"C1C2C1BE", x"BEC0C0BE",
									 -- x"C0BFBEBD", x"BDBEBFBF", x"C0BEBDBE", x"BFBFBFC0", x"C1C3C5C5", x"C4C3C5C8", x"C6C9CACA", x"CBCED0D0",
									 -- x"D3D1D2D6", x"D8D9DEE3", x"DEDFE0E0", x"DFDFE0E0", x"DCDEE0E0", x"DEDDDEE0", x"DEDEDDDC", x"DBDADADA",
									 -- x"D7D6D5D4", x"D4D2CFCD", x"CBCAC9C7", x"C3BFBDBC", x"BCB6B6B7", x"B4B1B0AD", x"A8AAABA8", x"A6A7A5A1",
									 -- x"A7A6A3A0", x"A0A09E9A", x"94939291", x"908F8D8B", x"89898682", x"81838481", x"807E807E", x"79777977",
									 -- x"73766F72", x"7270756F", x"6B696665", x"6463615E", x"5D5B5754", x"54565655", x"50525353", x"504E4F52",
									 -- x"51515151", x"504E5154", x"555B5455", x"575D575B", x"5B5E5F5F", x"62666561", x"63616261", x"5F626461",
									 -- x"66646160", x"61636464", x"63656460", x"60636361", x"5F606264", x"64626262", x"63626161", x"61616160",
									 -- x"6061615F", x"5E5E6062", x"5F5F6061", x"605F5D5D", x"5E5C5A57", x"56565859", x"55575652", x"4F4F5152",
									 -- x"54525150", x"504F5052", x"52535355", x"5556595C", x"5D60656A", x"6C6E7379", x"78797E7A", x"807F8787",
									 -- x"84817F81", x"83807C7A", x"77706D70", x"726E6967", x"67656465", x"625D5C5F", x"605C5859", x"5A5A5958",
									 -- x"55504C4D", x"4E4D4B4A", x"4A454142", x"4342403F", x"3E3C3B3A", x"3B393532", x"3537322D", x"30322F2D",
									 -- x"DBD9D5CF", x"CAC6C3C2", x"C3C3C4C4", x"C4C3C2C2", x"C1C4C7C7", x"C7C9CBCC", x"CECFD1D2", x"D3D2D1D1",
									 -- x"D2D1D0CF", x"CCC8C5C3", x"C4C3C4C4", x"BEB6B2B2", x"AFADABAA", x"AAA9A6A3", x"A7A4A2A3", x"A5A6A5A5",
									 -- x"A4A2A0A0", x"A1A2A1A0", x"9D999594", x"94929190", x"95969697", x"989A9D9E", x"9E9D9D9D", x"9FA1A2A2",
									 -- x"A2A4A5A7", x"A8AAABAC", x"AFAEADAE", x"AFB1B2B3", x"B7B9BBBD", x"BDBCBCBC", x"BEBFBFBE", x"BDBDBEBF",
									 -- x"C0BFBDBC", x"BBBBBABA", x"B9BCBEBD", x"BBBBBBBA", x"B6B4B3B2", x"B1B0AFAE", x"B1AFACAA", x"A9AAABAB",
									 -- x"A8A8A7A6", x"A5A5A6A7", x"A5A4A2A1", x"A09F9E9D", x"A09C9C9B", x"99999A98", x"97999997", x"95959595",
									 -- x"999A9B99", x"9A9C9E9E", x"9B9C9C9D", x"9E9FA0A1", x"9D9D9E9F", x"9F9F9F9F", x"9FA1A2A2", x"A2A19F9F",
									 -- x"9D9D9C9B", x"9B9B9D9E", x"9EA1A4A4", x"A5A8AAA9", x"ABACAEAF", x"AFB0B1B3", x"B2B4B7B8", x"B9BABBBD",
									 -- x"BFBEBEBF", x"C0C0BEBC", x"C2C1C0C0", x"C1C0BEBC", x"B9B7BABC", x"BBBDBFBE", x"BFBFBEBC", x"BDBFC2C2",
									 -- x"C2C1BFBE", x"BDBEBEBF", x"C1BFBDBE", x"BEBDBDBE", x"BFC0C0C1", x"C3C5C8C9", x"C5C6C7C9", x"CCD1D2D1",
									 -- x"D4D1D2D6", x"D8D9DDE2", x"DDDFE0E2", x"E1E1E0DF", x"DEDEDFDF", x"DFDFDEDE", x"DDDCDBD9", x"D8D7D7D7",
									 -- x"D3D3D3D3", x"D3D2CECB", x"C9C9C8C5", x"C1BFBDBC", x"BBB5B5B5", x"B2B0AEA9", x"A6A9A9A7", x"A6A7A5A1",
									 -- x"A6A4A2A2", x"9F9B9A9C", x"97979692", x"8D8A8A8A", x"8A8B8984", x"82848584", x"817E7F7E", x"79787874",
									 -- x"777B7375", x"75727770", x"706E6C6C", x"6B696562", x"5D5D5A56", x"54555656", x"50515150", x"4F4E4E4D",
									 -- x"504F5051", x"4F4E4F51", x"525A5658", x"585D5960", x"5C5D5C5C", x"6064625C", x"63616261", x"5E5F605B",
									 -- x"65625F5F", x"60626363", x"5E61615F", x"5F62615F", x"5D5F6161", x"62626261", x"5E5F5F5F", x"5E5D5D5D",
									 -- x"5E5E5D5C", x"5B5C5F62", x"5B5C5D5D", x"5C5B5958", x"5C5B5958", x"57565656", x"51535350", x"4F4F5151",
									 -- x"51505052", x"53535355", x"52535558", x"5856585B", x"5D60666B", x"6D6F757B", x"7E838B84", x"8581898B",
									 -- x"89858385", x"8684817E", x"7D767273", x"74706B68", x"6A666466", x"66636162", x"645F5A5A", x"5A585554",
									 -- x"56524E4D", x"4D4C4948", x"49494641", x"40403F3B", x"3D3B3938", x"39383634", x"3136332E", x"2F302F2F",
									 -- x"DBDAD8D3", x"CEC9C5C3", x"C3C3C3C4", x"C5C5C3C2", x"C2C4C6C6", x"C6C8C9C9", x"CBCDD0D2", x"D2D2D1D1",
									 -- x"D2D2D1D0", x"CECBC7C4", x"C7C6C4C3", x"BFB9B4B2", x"B1AEABAA", x"AAAAA7A5", x"A5A19FA0", x"A2A3A4A5",
									 -- x"A19F9D9C", x"9D9E9E9D", x"9D989594", x"94929190", x"95969696", x"97999C9C", x"9F9E9E9F", x"A0A0A09F",
									 -- x"A1A2A4A6", x"A7A8A9AA", x"AFAFAFAF", x"B0B2B3B4", x"B5B7B9BB", x"BCBBBBBB", x"BCBCBCBB", x"BBBDBFC0",
									 -- x"BFBDBBBA", x"BBBBBAB9", x"B7B9B9B8", x"B8B8B8B7", x"B6B4B1AF", x"AEAEADAD", x"ACABABAA", x"AAAAA9A8",
									 -- x"A8A7A6A4", x"A3A3A4A5", x"A3A3A2A1", x"A09F9D9C", x"9D9C9D9D", x"99999A98", x"94979997", x"95959798",
									 -- x"96999A9A", x"9A9B9B9A", x"97989A9A", x"9A9B9D9E", x"9D9D9E9E", x"9E9E9FA0", x"9F9FA0A1", x"A1A09F9E",
									 -- x"9B9B9B9B", x"9B9B9B9C", x"9DA0A2A1", x"A3A7A9A8", x"AAAAACAE", x"AEAEAFB0", x"B1B3B5B7", x"B9BABBBB",
									 -- x"BABABBBC", x"BDBDBBBA", x"BFBEBDBD", x"BCBAB8B8", x"B9B7B9BA", x"B8BABCBA", x"BBBBBBBA", x"BBBEC1C3",
									 -- x"C3C2C0BF", x"BEBDBDBE", x"C1BEBDBE", x"BEBEBEBF", x"BFBFBFC0", x"C2C6C9C9", x"C6C6C7C9", x"CDD2D3D2",
									 -- x"D1D2D4D7", x"D9DADCDE", x"DDDEE0E1", x"E2E1E0DF", x"E0DFDEDE", x"DFDFDEDC", x"DDDCDAD8", x"D6D5D4D4",
									 -- x"D1D1D1D1", x"D2D0CDCA", x"C5C6C5C2", x"BFBEBDBC", x"B9B4B2B2", x"AFAEABA6", x"A6A7A8A7", x"A6A6A5A3",
									 -- x"A5A2A2A2", x"9F9A999C", x"98989792", x"8C898A8C", x"8B8D8C87", x"84868785", x"817D7C7C", x"78777672",
									 -- x"767A787A", x"79777671", x"75727070", x"6F6B6663", x"5D5E5C57", x"54545555", x"4F504F4E", x"4F4F4D4B",
									 -- x"514C4A4C", x"50504D4C", x"4A52545A", x"585B595D", x"5C5C5B5B", x"5E605E5B", x"605F6060", x"5D5F5F5B",
									 -- x"5F5E5D5D", x"5F616161", x"5B5D5F5F", x"5F605E5C", x"5B5C5D5D", x"5D5E5F5E", x"5A5A5C5D", x"5C59595A",
									 -- x"59595959", x"5A5B5B5C", x"5B5B5957", x"57595958", x"5B5A5857", x"56555352", x"504F4C4D", x"5154534F",
									 -- x"4F4F5052", x"52515152", x"5254585C", x"5B575659", x"5F616469", x"6C70767B", x"84888D8A", x"8B8B8F8E",
									 -- x"8D898787", x"87848280", x"837F7A76", x"74726E6B", x"6B686769", x"6A686461", x"605D5C5C", x"5C595553",
									 -- x"5753504F", x"4D4A4746", x"46494741", x"3F41403C", x"3B393737", x"37383736", x"2F35332F", x"2F2F2E30",
									 -- x"DCDDDCD8", x"D3CDC8C6", x"C5C4C3C3", x"C4C5C5C4", x"C4C5C5C5", x"C7CAC9C7", x"CACDD0D1", x"D2D1D2D2",
									 -- x"D3D3D3D3", x"D2CFCBC8", x"C8C7C4C2", x"C1BFBBB6", x"B4B0ABA9", x"A9A9A7A5", x"A29F9D9E", x"9F9FA0A2",
									 -- x"9C9B9998", x"999A9B9B", x"9B969393", x"94939393", x"94969897", x"989A9B9B", x"9E9FA0A1", x"A1A09F9E",
									 -- x"A0A2A4A5", x"A6A7A8A9", x"ADAEAFB0", x"B0B1B3B4", x"B3B4B6B8", x"B9B9BABB", x"B9B9B9BA", x"BABCBEBF",
									 -- x"BFBCBAB9", x"BABBBAB8", x"B7B7B7B5", x"B6B8B8B6", x"B6B4B0AD", x"ACACACAB", x"AAA9A9A9", x"A9A8A7A6",
									 -- x"A7A7A6A5", x"A3A2A3A3", x"A1A1A1A1", x"A1A09E9D", x"9B9B9E9E", x"98979998", x"95979896", x"95979899",
									 -- x"95989A99", x"999A9A98", x"97979797", x"999A9B9C", x"9C9D9D9C", x"9C9C9EA0", x"9E9E9E9E", x"9F9E9E9D",
									 -- x"9A9B9B9B", x"9B9C9D9E", x"9F9FA0A2", x"A3A4A6A8", x"A9A8A8AB", x"ADADAEB0", x"B2B1B1B3", x"B6B8B8B8",
									 -- x"B5B6B8B9", x"B9B8B7B7", x"BBB9B8B8", x"B7B5B6B8", x"BCB9B9B9", x"B6B6B8B6", x"BABABBBB", x"BBBCBFC1",
									 -- x"C1C0C0BF", x"BFBEBFBF", x"C1BFBDBE", x"BFBFBFC1", x"C0C3C3C2", x"C2C5C7C7", x"C6C7C8C9", x"CBCFD1D0",
									 -- x"CFD1D4D5", x"D7DADCDC", x"DEDEDFE0", x"E1E1E1E0", x"DFDFDFDE", x"DEDDDCDB", x"DBDAD9D7", x"D5D4D3D2",
									 -- x"D1D0CFCF", x"CFCDCBC8", x"C5C6C4C0", x"BEBEBEBC", x"B9B3B0AF", x"ADADACA6", x"A8A7A7A8", x"A8A6A5A6",
									 -- x"A4A4A3A1", x"9F9D9B99", x"96969592", x"8E8C8D8E", x"8B8C8B87", x"86878682", x"7F7C7C7B", x"78777773",
									 -- x"75777C7B", x"7A7B7776", x"79757272", x"716D6867", x"6162605C", x"58585756", x"52535351", x"51514F4C",
									 -- x"514C494B", x"4E4F4E4C", x"4A4E5159", x"54585657", x"5A59595B", x"5A595A5C", x"5E5D5E5D", x"5C5F605D",
									 -- x"5B5B5C5E", x"5F5F5E5E", x"5A5A5C5E", x"5E5C5A5A", x"5B5C5C5A", x"595B5C5C", x"5857585B", x"5C5A5858",
									 -- x"57565657", x"58595857", x"59595654", x"54565755", x"57565554", x"54535251", x"504D4B4B", x"5054534F",
									 -- x"4F4E4F51", x"52504F50", x"5555595D", x"5C595A5F", x"64636468", x"6D73797E", x"868B8C8E", x"8E949391",
									 -- x"918E8B8A", x"89878586", x"86858079", x"75757472", x"6D6D6C6B", x"6A686561", x"5E5C5B5C", x"5C5A5959",
									 -- x"57545250", x"4E494645", x"45444241", x"4141403D", x"39383837", x"36363535", x"30333230", x"312F2D2E",
									 -- x"DFE0DFDC", x"D6D0CCCA", x"C7C5C3C3", x"C4C5C6C6", x"C5C6C5C5", x"C8CBCAC7", x"CBCDD0D1", x"D2D2D3D4",
									 -- x"D4D4D4D5", x"D4D2CECB", x"C6C6C4C2", x"C3C5C1BB", x"B6B1ABA8", x"A8A8A6A4", x"A29F9D9E", x"9E9C9D9F",
									 -- x"9B9A9898", x"999A9B9C", x"99959292", x"94949495", x"90949797", x"989A9A99", x"9D9FA1A2", x"A1A09E9E",
									 -- x"A0A2A4A5", x"A6A7A8A8", x"AAACAEAF", x"AEAFB1B3", x"B2B3B4B5", x"B6B7BABB", x"B7B8B9B9", x"B9BABCBD",
									 -- x"C0BDB9B8", x"BABAB9B8", x"B9B9B7B6", x"B7B9B9B7", x"B7B4B0AC", x"ABAAABAB", x"ABA9A7A6", x"A5A6A6A6",
									 -- x"A4A5A5A4", x"A2A0A0A0", x"9E9E9FA0", x"A09F9D9C", x"9A9B9E9D", x"97969999", x"9D9C9A97", x"96969594",
									 -- x"96989998", x"98999A99", x"9B999799", x"9C9E9E9D", x"9C9C9C9B", x"9A9A9C9E", x"9F9E9C9C", x"9C9D9D9E",
									 -- x"9B9B9C9C", x"9D9EA0A1", x"A49F9FA4", x"A5A1A3A9", x"A9A6A6A9", x"ACADAFB2", x"B3B1AEB0", x"B3B6B6B5",
									 -- x"B5B7B9B9", x"B8B6B5B5", x"B7B6B5B5", x"B5B5B8BD", x"B9B6B6B6", x"B3B4B6B4", x"BABBBCBD", x"BDBCBEC0",
									 -- x"BDBEBEBF", x"C0C0C1C1", x"C3C0BEBF", x"BFBFC0C1", x"C2C6C8C5", x"C3C3C5C5", x"C5C8C9C9", x"C9CBCDCE",
									 -- x"CED1D2D0", x"D2D8DCDB", x"DFDFDEDF", x"E0E1E2E2", x"DEDFE0DF", x"DCDBDBDB", x"D9D9D8D7", x"D6D4D4D3",
									 -- x"D3D1CECD", x"CCCBC9C8", x"C7C8C6C1", x"BEBEBEBC", x"BAB4B0AE", x"ADAEAEA9", x"A9A7A7A9", x"A9A6A6A9",
									 -- x"A3A6A49F", x"9FA29E97", x"98979592", x"908E8D8C", x"8A8A8885", x"8687847E", x"7F7D7D7D", x"78787977",
									 -- x"79777F7A", x"787C7578", x"7D797676", x"75716E6E", x"67666460", x"5F5E5B58", x"55575754", x"52514F4C",
									 -- x"504E4D4D", x"4C4C4E51", x"52505259", x"52575654", x"5656585A", x"5754575E", x"5E5C5C5C", x"5A5E615E",
									 -- x"5B5C5E5F", x"5F5D5C5A", x"5B595A5D", x"5D595859", x"5D5E5D59", x"585B5C5C", x"5956565A", x"5D5C5A59",
									 -- x"59565354", x"56585756", x"54555452", x"5253524E", x"53515051", x"52525251", x"4E4F4E4C", x"4C4F5151",
									 -- x"4E4E5053", x"54545456", x"5957595C", x"5C5C6168", x"69656469", x"70777D82", x"8A918F93", x"8E969392",
									 -- x"95939190", x"8E8C8D8E", x"8587847A", x"76797A78", x"71727069", x"66666562", x"64605D5B", x"59585A5D",
									 -- x"56545351", x"4E494645", x"48423E41", x"423E3A39", x"39393938", x"36343232", x"32333030", x"322F2B2D",
									 -- x"E1E2E2DE", x"D9D5CFCA", x"C8C6C5C4", x"C4C3C5C7", x"C7C6C6C7", x"C8C7C7C8", x"CDCDCDCF", x"D1D2D3D3",
									 -- x"D7D7D6D4", x"D3D1CECA", x"CAC5C1C0", x"C2C2C0BD", x"B7B3ADA7", x"A8AAA8A2", x"A1A09D9B", x"9A9A9B9D",
									 -- x"9A999897", x"98999895", x"95969392", x"94939398", x"91929294", x"989C9B97", x"9D9E9FA0", x"9F9F9E9E",
									 -- x"9EA0A3A5", x"A6A8A9AA", x"AAAAABAD", x"AFB0AFAD", x"B1B2B3B4", x"B5B7BABC", x"B7B7B7B7", x"B8BABDBF",
									 -- x"BEBEBCB9", x"BABBBAB7", x"B8B9B9B9", x"B8B7B8B9", x"B6B1AEAB", x"AAACABA4", x"A5A8A6A1", x"A1A5A5A0",
									 -- x"A3A3A2A0", x"9F9E9FA0", x"9FA0A09F", x"9E9D9D9D", x"9C9C9C9B", x"9A999A9A", x"999A9A99", x"97959596",
									 -- x"999B9B99", x"99999794", x"989B9D9C", x"9A999B9E", x"9D9D9997", x"999A9B9F", x"9B99999B", x"9C9C9C9D",
									 -- x"9D9D9C9E", x"9FA09F9E", x"9FA0A1A1", x"A2A3A4A5", x"A4A5A7A9", x"ABADAEAE", x"B2B2B2B0", x"AFAFB1B4",
									 -- x"B0B2B4B6", x"B6B6B6B6", x"B7B5B5B4", x"B2B6B8B4", x"B6B5B5B4", x"B6B7B6B3", x"B3B5B6B8", x"B9BBBFC2",
									 -- x"C0C1C2C3", x"C1C0C1C4", x"C2C1C0BF", x"BEBFC0C2", x"C4C7C4C3", x"C6C3BFC3", x"C5C5C6C8", x"C9C9CCCF",
									 -- x"D0D1D2D2", x"D3D3D5D7", x"D5D9DDE1", x"E2E1DFDE", x"DFDFDFDE", x"DBD9D9D9", x"D7D5D4D3", x"D4D4D1CF",
									 -- x"CFCFCECB", x"C9C7C6C4", x"C7C6C3BF", x"BCBCBCBC", x"B8B5B1AF", x"AFAFAEAD", x"A8A6A6A9", x"A9A5A4A7",
									 -- x"A3A4A29E", x"9EA1A09C", x"9B9A9795", x"92908F8F", x"89888788", x"86828082", x"807E7B79", x"797B7D7F",
									 -- x"7C7F7C79", x"7D7E7A78", x"7B7B7980", x"77736D72", x"6E696565", x"64605C5A", x"55565553", x"51504F4F",
									 -- x"544B474B", x"4E4B4C50", x"4F4B5056", x"5350545A", x"5657565A", x"5858605E", x"5D5D5C59", x"595A5C5B",
									 -- x"585E625F", x"5A5A5B5D", x"58595C5D", x"5A57575A", x"595B5D5C", x"5B595959", x"59575656", x"59595754",
									 -- x"52525253", x"53535251", x"57535153", x"524D4A4A", x"4C4D4F4E", x"4C4C4D4E", x"4B4D4E4F", x"50505050",
									 -- x"51535557", x"5757585A", x"5C615F5D", x"646A6864", x"67696B6C", x"6E75818A", x"93989994", x"93989A98",
									 -- x"99989592", x"91918F8B", x"8885827F", x"7E84847B", x"76706F6A", x"696A6464", x"6261605E", x"5D5B5B5A",
									 -- x"5558514E", x"514D4648", x"4744403E", x"3F3E3C3A", x"38383634", x"33343433", x"2F2E2F30", x"32312E2B",
									 -- x"E2E3E3E1", x"DDD9D2CC", x"CCC9C6C4", x"C3C3C6CA", x"C3C3C4C6", x"C6C6C7C9", x"CCCDCFD1", x"D2D3D4D5",
									 -- x"D5D6D5D4", x"D4D3CEC9", x"C8C5C1C1", x"C2C1BFBC", x"B7B3ADA9", x"A9AAA8A5", x"A19F9C9B", x"9C9D9D9C",
									 -- x"97989896", x"96969694", x"94959291", x"928F8E92", x"91929292", x"94979693", x"98999A9B", x"9C9D9D9E",
									 -- x"9E9FA0A1", x"A2A3A5A6", x"A8A8A9AB", x"ADAFAFAF", x"B1B1B3B4", x"B6B7B8B9", x"B7B7B7B7", x"B7B8BBBD",
									 -- x"BEBEBDBB", x"BBBBBAB8", x"B8B8B9B8", x"B7B6B7B7", x"B6B1AFAB", x"A9ABABA5", x"A6A7A5A1", x"A1A3A29E",
									 -- x"9FA09F9F", x"9E9FA0A1", x"9FA0A0A0", x"9F9E9E9E", x"9C9C9C9B", x"9A999999", x"98999998", x"97969797",
									 -- x"9A9B9A99", x"99999895", x"979A9C9C", x"9A999A9C", x"9C9D9A99", x"9B9B9B9E", x"9B99999B", x"9C9C9B9C",
									 -- x"9D9C9C9C", x"9E9FA09F", x"9FA0A2A2", x"A2A3A3A4", x"A4A5A7A8", x"AAACADAD", x"B5B4B2B1", x"B1B1B2B2",
									 -- x"B1B1B0B0", x"B0B1B3B5", x"B4B2B2B2", x"B0B4B6B2", x"B3B5B6B8", x"B9B9B5B0", x"B4B5B5B6", x"B7BABEC1",
									 -- x"C1C0C2C3", x"C3C3C5C8", x"C7C5C2C1", x"C1C3C5C7", x"C5C5C3C3", x"C5C2C1C3", x"C8C7C8CA", x"CACACCCF",
									 -- x"D0D1D2D3", x"D2D2D3D4", x"D8D9DBDC", x"DCDDDDDE", x"DEDEDCDA", x"D8D8D9DA", x"D7D5D3D3", x"D3D2D0CE",
									 -- x"C9C9C9C9", x"C8C8C8C8", x"C3C3C2C0", x"BDBBB9B8", x"B8B6B3B1", x"B1B0AEAC", x"A8A5A4A7", x"A7A4A5A8",
									 -- x"A3A2A09D", x"9C9C9A98", x"9B989593", x"918E8A88", x"8F8C8A88", x"85828182", x"817E7C7B", x"7B7B7C7C",
									 -- x"807E7C7F", x"817C7C85", x"827D7C7C", x"7D787675", x"736E6866", x"635F5C5C", x"56565655", x"53525252",
									 -- x"504F4D4D", x"4D4C4B4A", x"4A494D51", x"50505251", x"50535559", x"57555B58", x"5A595B5D", x"5C595A5E",
									 -- x"605E5C5B", x"5E615E5A", x"5A5B5C5D", x"5B575759", x"57575758", x"58575655", x"59575655", x"5554524F",
									 -- x"51504F50", x"5151504F", x"4F4B4B4D", x"4D4A4849", x"494B4D4D", x"4B494949", x"4E4E4F52", x"54555452",
									 -- x"5557595A", x"595A5B5C", x"60616063", x"6A6B696C", x"6D6F7071", x"73798289", x"8B949C9D", x"9B9B9997",
									 -- x"9B9B9994", x"918F8E8C", x"89868582", x"8083837D", x"7A75746E", x"6B6A6363", x"6564615E", x"5C595756",
									 -- x"5557514E", x"514E4849", x"4744413F", x"3F3E3C3A", x"37363331", x"3234322F", x"302F2E2E", x"2E2E2C2B",
									 -- x"E3E4E4E3", x"E1DDD5CE", x"CDC9C7C5", x"C5C5C7CA", x"C4C4C5C6", x"C6C5C7CA", x"CACDD0D1", x"D2D3D5D7",
									 -- x"D5D6D5D5", x"D5D3CEC8", x"C6C4C2C1", x"C0BFBDBB", x"BAB5AFAD", x"ABAAAAAA", x"A4A09D9D", x"9FA09E9C",
									 -- x"97999A97", x"96959595", x"94959493", x"938F8C8F", x"91929291", x"91929291", x"94959697", x"989A9B9D",
									 -- x"9E9F9FA0", x"A1A3A5A6", x"A6A7A8AA", x"ABACAEAF", x"AFAFB0B3", x"B4B5B5B5", x"B6B7B8B8", x"B6B6B9BB",
									 -- x"BCBDBEBC", x"BBBAB9B8", x"B7B8B8B8", x"B7B7B7B7", x"B6B2B0AD", x"A9ABABA8", x"A6A5A3A2", x"A2A09F9E",
									 -- x"9E9E9E9E", x"9E9FA0A1", x"9F9FA0A1", x"A0A09F9E", x"9D9D9D9D", x"9C9A9998", x"999A9A9A", x"9A9A9B9C",
									 -- x"9A9A9A98", x"99999896", x"96989A9B", x"9A9A9999", x"9B9D9C9B", x"9D9C9B9D", x"9B99999B", x"9C9B9B9C",
									 -- x"9D9C9B9C", x"9D9FA0A0", x"9EA0A2A3", x"A3A4A4A4", x"A5A5A7A8", x"A9ABACAC", x"B3B1AFAF", x"B1B1B0AF",
									 -- x"B0B0AFAF", x"AFB0B2B4", x"B1AFB0B0", x"AFB2B4B1", x"B0B2B4B6", x"B7B6B2AD", x"B4B4B4B3", x"B4B7BCBF",
									 -- x"C2C1C1C3", x"C4C5C7C9", x"C9C7C5C5", x"C7C9CBCB", x"CAC6C6C7", x"C5C5C7C7", x"C8C7C6C8", x"CACACACC",
									 -- x"D0D1D2D2", x"D2D1D2D2", x"D8D8D8D8", x"D8D9DADB", x"DBDBDAD9", x"D7D7D8D9", x"D6D4D3D2", x"D2D1CFCD",
									 -- x"CAC9C8C8", x"C7C7C7C7", x"C1C0C0BF", x"BDB9B7B5", x"B6B5B3B2", x"B1B0AEAC", x"A6A4A5A8", x"A8A6A6A8",
									 -- x"A5A2A09E", x"9C9A9898", x"97959392", x"93928D89", x"8E8C8987", x"84818080", x"82817E7D", x"7D7D7C7C",
									 -- x"807F7F81", x"827E828E", x"89818079", x"817C7D77", x"76736E6A", x"65605D5C", x"57575756", x"55545454",
									 -- x"50545450", x"4E4F4E4B", x"494A4E4F", x"4F52524B", x"5054555A", x"57545A56", x"58575A5E", x"5C585A61",
									 -- x"61626160", x"6060605E", x"5C5B5B5C", x"5B585758", x"56555454", x"56565452", x"59595856", x"54524F4E",
									 -- x"514F4D4E", x"50515150", x"4E4C4C4F", x"4F4D4D4E", x"4D4E5050", x"504F4E4E", x"51515255", x"595B5957",
									 -- x"5B5D5E5F", x"5F5F6162", x"6662626A", x"716D6D75", x"74757575", x"777C8389", x"8A929DA1", x"A09D9C9C",
									 -- x"9E9E9C97", x"9391908F", x"8D898887", x"8383827E", x"7B777670", x"6C6A6363", x"63615F5D", x"5B5A5958",
									 -- x"5556514F", x"504E494A", x"4644413F", x"3D3C3A39", x"37353230", x"3133312D", x"31302E2D", x"2C2C2C2D",
									 -- x"E6E6E5E4", x"E3DFD7CF", x"CBC9C7C8", x"C8C7C7C8", x"C6C6C6C7", x"C5C3C5C8", x"C7CBCECE", x"CECFD4D8",
									 -- x"D8D7D6D4", x"D5D4CEC8", x"C5C4C2BF", x"BEBCBCBB", x"BCB7B3B2", x"AFABABAD", x"A8A5A1A0", x"A1A19F9D",
									 -- x"9B9C9C9A", x"99999896", x"93949393", x"94918E91", x"91939493", x"92919191", x"92939596", x"9697999A",
									 -- x"9C9D9FA0", x"A2A4A6A7", x"A5A7A9AA", x"AAAAABAC", x"AFAFB0B2", x"B4B5B5B4", x"B5B7B9B8", x"B7B6B8BB",
									 -- x"B9BBBDBD", x"BBBAB9B9", x"B8B8B8B8", x"B8B8B8B8", x"B5B2B2B1", x"ACABACAA", x"A6A3A2A4", x"A3A09E9F",
									 -- x"A0A0A0A0", x"9F9FA0A0", x"9F9FA0A1", x"A1A1A09F", x"9F9F9F9F", x"9E9C9997", x"9A9A9A9A", x"9B9B9C9D",
									 -- x"9A999898", x"98999898", x"9898999A", x"9A9A9998", x"9B9D9C9B", x"9E9D9C9E", x"9B9A999B", x"9C9B9B9C",
									 -- x"9D9D9C9C", x"9D9E9E9F", x"9D9FA1A3", x"A4A5A7A8", x"A5A6A7A8", x"A9AAACAC", x"ADADADAE", x"AFB0B0AF",
									 -- x"ACADAFB0", x"B1B0B1B1", x"B0AEAFB0", x"AFB1B3B1", x"B1B2B2B1", x"B1B2B0AE", x"B2B2B2B2", x"B3B5BABD",
									 -- x"C3C1C1C4", x"C6C6C7C8", x"CAC8C7C9", x"CCCECECD", x"CEC7C9CA", x"C5C6CBC9", x"C8C5C4C7", x"C9C9CACA",
									 -- x"D0D0D0D0", x"D0D1D2D2", x"D4D5D7D7", x"D7D7D7D7", x"D7D8D9DA", x"D9D8D6D5", x"D4D3D2D1", x"D1D0CECD",
									 -- x"CBC9C7C6", x"C5C3C2C3", x"C2BFBDBC", x"BAB8B6B6", x"B3B2B0AF", x"AFAEACAB", x"A6A6A8AB", x"ABA8A6A6",
									 -- x"A8A4A1A1", x"9F9B9A9C", x"97969595", x"9696938F", x"8A898887", x"8683807E", x"81807F7E", x"7D7D7E7E",
									 -- x"7C828380", x"83878A8D", x"8C86827C", x"807E7C74", x"74747370", x"6A635E5C", x"59585858", x"56545455",
									 -- x"52545350", x"4F505151", x"4F4F5253", x"5253534D", x"56565558", x"57565C57", x"5A595B5D", x"5C5A5D62",
									 -- x"61656866", x"63606060", x"5A595859", x"5A595857", x"57565555", x"56555452", x"56575857", x"54525050",
									 -- x"504D4B4C", x"4F515150", x"4C4B4B4D", x"4D4C4C4D", x"4D4D4E4F", x"50525354", x"5455565A", x"5D5F605F",
									 -- x"60616364", x"64656869", x"6A67666E", x"7471727B", x"7D7D7C7B", x"7B7F878D", x"9093999E", x"9E9C9FA3",
									 -- x"9F9E9D9B", x"98969492", x"908A8889", x"8684817C", x"7A75746E", x"6A696364", x"615F5D5B", x"5B5B5A59",
									 -- x"5655524F", x"4F4C4A49", x"4443413E", x"3B393837", x"37363331", x"3132302D", x"2F2F2D2B", x"2A2A2C2D",
									 -- x"E7E7E5E4", x"E3E1DBD5", x"CFCCCACA", x"C9C7C6C6", x"C6C5C4C4", x"C3C1C2C4", x"C4C7C9C9", x"C8CAD0D5",
									 -- x"D8D7D5D4", x"D4D4D1CC", x"C6C5C2BE", x"BCBBBBBB", x"BCB8B6B5", x"B2ACAAAC", x"A9A7A4A1", x"A0A0A1A2",
									 -- x"A09F9D9C", x"9D9E9A96", x"93949392", x"94918F92", x"95969899", x"96939293", x"91929495", x"95969797",
									 -- x"9A9B9EA0", x"A1A3A4A5", x"A3A6A9AA", x"AAA9AAAB", x"B1B1B1B2", x"B4B5B6B6", x"B5B7B9B9", x"B8B8BABC",
									 -- x"B9BBBDBE", x"BDBCBCBD", x"BABAB9B8", x"B8B7B6B6", x"B3B1B2B2", x"ADABACA9", x"A8A4A3A5", x"A4A09E9F",
									 -- x"A1A1A1A0", x"9F9F9F9F", x"9F9F9FA0", x"A1A1A09F", x"A0A0A0A0", x"A09E9B98", x"99999999", x"99999999",
									 -- x"99989797", x"98989899", x"99999899", x"9A9A9999", x"9B9D9B9B", x"9D9E9DA0", x"9C9A9A9C", x"9D9C9B9C",
									 -- x"9D9D9D9D", x"9D9C9C9C", x"9FA0A1A2", x"A3A5A8AA", x"A6A6A7A8", x"A9AAACAC", x"AAACAEAF", x"AFAFB0B1",
									 -- x"AAABAEAF", x"AFAEADAD", x"B0ADAFB0", x"ADAFB1B0", x"B2B2B1AF", x"AEB0B0AF", x"AFB0B1B2", x"B3B5B8BB",
									 -- x"C1C0C1C6", x"C9CACBCC", x"CDCBC9CB", x"CED1D2D1", x"CEC8C9CA", x"C5C6CAC8", x"C9C7C6C8", x"C9C9C9CA",
									 -- x"CECDCDCD", x"CED0D2D3", x"D2D3D4D5", x"D5D5D6D6", x"D6D7D8D9", x"D9D7D4D3", x"D2D1D0D0", x"D0CFCECD",
									 -- x"C7C5C3C3", x"C2C1C1C3", x"C1BEBCBC", x"BAB7B5B5", x"B1B0AEAC", x"ACACACAC", x"A8A8A9AA", x"AAA7A5A5",
									 -- x"A8A4A2A2", x"9F9B9A9C", x"999A9996", x"94949391", x"8B8A8887", x"86848280", x"7D7E7E7C", x"7B7C7F83",
									 -- x"7D828383", x"898C8B8B", x"8D8B8382", x"7D7E7671", x"73747571", x"6B65615E", x"5B595858", x"56535254",
									 -- x"53504F50", x"51505052", x"55525456", x"52515252", x"59565357", x"58585C56", x"5A5E5F60", x"62646461",
									 -- x"68666463", x"63625F5D", x"59585656", x"58585756", x"56575857", x"55535353", x"52545555", x"53525353",
									 -- x"4E4C4A4A", x"4C4D4D4C", x"4C4B4B4C", x"4D4C4D4E", x"4D4F5254", x"56575859", x"585A5D5F", x"61646769",
									 -- x"65666767", x"68696C6E", x"6E6E6D70", x"75767980", x"83868785", x"8384898E", x"9392959A", x"9C9C9EA2",
									 -- x"9F9D9B9B", x"9B999491", x"91898889", x"8886827C", x"7A74726B", x"67686365", x"64615E5B", x"5A585655",
									 -- x"5653514F", x"4C4A4947", x"4443413E", x"3B383736", x"35363532", x"3030302E", x"2C2C2B2A", x"29292A2B",
									 -- x"E8E8E7E5", x"E5E4E0DB", x"D7D2CDCA", x"C8C7C6C7", x"C6C4C3C3", x"C3C2C3C5", x"C2C4C6C5", x"C4C6CCD0",
									 -- x"D5D5D4D3", x"D4D5D4D1", x"CBC8C4C0", x"BDBCBCBD", x"BAB8B7B5", x"B2ADAAA9", x"A7A6A4A2", x"A1A1A3A5",
									 -- x"A3A19E9E", x"A0A09C96", x"97989695", x"96939296", x"9B9B9C9D", x"9A969495", x"91929394", x"94959697",
									 -- x"9B9C9FA0", x"A1A2A3A3", x"A2A4A6A8", x"A9AAAAAB", x"ADAEAFB0", x"B1B2B4B5", x"B5B6B7B9", x"BABBBDBE",
									 -- x"BDBDBDBF", x"BFBEBFC0", x"BEBCBAB9", x"B7B6B4B2", x"B1AFB0B1", x"ACAAAAA9", x"ABA7A5A5", x"A4A09E9F",
									 -- x"A0A0A0A0", x"9F9E9F9F", x"9F9E9E9E", x"A0A09F9E", x"A0A0A0A0", x"A19F9C9A", x"9B9A9A9A", x"9A9A9998",
									 -- x"99979798", x"9998999A", x"9A999999", x"999A9A99", x"9C9D9B9A", x"9D9D9DA0", x"9D9B9B9C", x"9D9C9C9D",
									 -- x"9C9D9E9D", x"9C9B9B9B", x"A0A1A1A1", x"A2A4A6A9", x"A6A6A6A7", x"A8A9AAAB", x"A8AAACAC", x"ABABADAE",
									 -- x"AEAEAEAD", x"ACADAEAF", x"B0ACADAE", x"ABABAEAE", x"ADAFAFAE", x"ADAEADAC", x"ADAEB0B1", x"B3B5B9BC",
									 -- x"BDBEC1C6", x"CBCDD1D3", x"D2CFCBCA", x"CCD0D3D4", x"CFCBCACA", x"C7C6C7C7", x"C8C6C5C6", x"C7C6C7C8",
									 -- x"CBCAC9CA", x"CCCED0D1", x"D1D1D1D1", x"D1D3D5D7", x"D7D6D5D4", x"D4D4D3D2", x"CFCFCFCE", x"CDCCCBCB",
									 -- x"C8C5C3C4", x"C3C0C0C2", x"BEBBBABC", x"BBB6B2B1", x"B0AFADAB", x"AAAAABAB", x"A9A8A7A6", x"A5A4A3A4",
									 -- x"A5A3A19F", x"9C999899", x"95979692", x"91939392", x"8E8C8884", x"83838280", x"7E7E7E7D", x"7C7E8388",
									 -- x"82808188", x"8D89868C", x"8E8D8486", x"7C7C7270", x"7475746F", x"6A666462", x"5D5A595A", x"57535254",
									 -- x"54515155", x"56535152", x"58535456", x"52505355", x"5958565B", x"5D5D5F58", x"5B626667", x"6A6E6A61",
									 -- x"67656360", x"5D5B5C60", x"5B5A5856", x"56575755", x"55575958", x"55535252", x"52545555", x"55545557",
									 -- x"4F4F4E4D", x"4D4D4C4B", x"4D4E4E4F", x"4F505153", x"51555B5E", x"5E5D5C5C", x"5E616567", x"686A6E72",
									 -- x"6C6D6D6C", x"6C6D6F71", x"73777776", x"7A7E8185", x"888B8F8F", x"8C8A8A8B", x"9090949B", x"9E9C9A9B",
									 -- x"A09C999A", x"9B97918D", x"8F8A8889", x"8787837C", x"7B747069", x"67686364", x"64615C59", x"58575452",
									 -- x"5551504E", x"48474744", x"4442403D", x"3B393735", x"31343431", x"2E2E2E2E", x"2C2C2C2C", x"2C2B2B2A",
									 -- x"E9E9E8E6", x"E4E3E0DC", x"DAD4CECA", x"C9C7C7C8", x"C7C3C1C3", x"C4C4C4C5", x"C2C4C5C5", x"C4C5C9CC",
									 -- x"D0D3D4D3", x"D3D4D4D3", x"D0CCC8C4", x"C1C0BFBE", x"BABAB8B5", x"B2B0ACA9", x"A9A7A4A3", x"A4A5A6A6",
									 -- x"A4A3A1A0", x"A1A19D98", x"9B9C9A9A", x"9B979699", x"9F9D9D9D", x"9B989798", x"96969594", x"94949698",
									 -- x"9B9C9E9F", x"A0A1A2A3", x"A3A3A3A5", x"A7A9AAAA", x"A8ABAEB0", x"AFAFB1B4", x"B5B5B5B7", x"BABDBEBE",
									 -- x"C0BEBDBE", x"BFBEBFC1", x"C0BFBCBA", x"B9B7B5B3", x"B3AFAFB0", x"ACABABAA", x"AAA8A6A5", x"A3A2A1A0",
									 -- x"A0A1A1A1", x"A09F9F9F", x"A09E9C9D", x"9E9F9E9D", x"9F9F9E9F", x"A0A09D9B", x"9D9D9C9D", x"9D9D9A99",
									 -- x"99979799", x"9A9A9A9B", x"99999A9A", x"9A999999", x"9C9E9C9A", x"9D9D9C9E", x"9E9C9C9D", x"9E9D9D9D",
									 -- x"9D9D9D9D", x"9B9B9B9C", x"9F9FA0A0", x"A1A2A5A6", x"A7A7A6A6", x"A6A7A8A8", x"A6A7A8A8", x"A9AAABAC",
									 -- x"AEAEADAC", x"ACADB0B2", x"B1ADADAD", x"A8A8ABAD", x"A8AAACAB", x"ABACACAB", x"ACADAFB0", x"B2B6BABE",
									 -- x"BEBEC1C5", x"C8CBD0D5", x"D3D1CECB", x"CBCDCFD1", x"CFCFCCCB", x"CAC6C4C6", x"C4C3C3C5", x"C5C4C6C8",
									 -- x"C8C7C7C8", x"CACBCBCB", x"CFCFD0D0", x"D0D1D2D4", x"D4D3D1D1", x"D1D1D0CF", x"CECECDCC", x"CAC8C7C7",
									 -- x"C9C5C4C5", x"C3BEBDBF", x"BCB8B7B9", x"B9B3AFAF", x"AEADACAA", x"A8A7A7A8", x"A7A7A6A4", x"A3A2A1A0",
									 -- x"A2A3A19D", x"9A999898", x"9294928F", x"90949491", x"8D8C8985", x"8484817D", x"807F7D7C", x"7E818587",
									 -- x"80818387", x"8781828C", x"918A8382", x"7E797473", x"7576746F", x"6A686562", x"5F5C5B5C", x"59545355",
									 -- x"54565857", x"57575656", x"5D595857", x"55585B59", x"5C5C5B60", x"60606560", x"60656A6C", x"6D6E6964",
									 -- x"63636461", x"5B575B61", x"5C5C5A57", x"57585857", x"57585A5B", x"5A585654", x"57575656", x"55555656",
									 -- x"4F505252", x"504F4F4F", x"4E4F5050", x"50515354", x"52585E60", x"5E5C5C5E", x"64676C6F", x"71737678",
									 -- x"75757473", x"72737678", x"797F8182", x"8587898D", x"8F919395", x"9594918F", x"9194989B", x"9D9C9C9C",
									 -- x"A29D9A9A", x"9994908D", x"8E8D8D8A", x"8585837B", x"7A726E68", x"67696363", x"605C5856", x"56565452",
									 -- x"524D4E4C", x"45444642", x"42403D3B", x"3A393533", x"30323230", x"2E2E2D2C", x"2D2C2B2C", x"2C2C2A29",
									 -- x"E9EAEAE6", x"E3E0DDDA", x"D7D2CDCB", x"CAC8C7C6", x"C6C2BFC1", x"C3C3C3C3", x"C2C4C6C6", x"C6C6C8CA",
									 -- x"CED2D4D4", x"D3D3D3D2", x"D3D0CBC8", x"C6C4C1BF", x"BBBCB9B4", x"B3B3B0AA", x"ACA9A6A6", x"A8A9A7A5",
									 -- x"A5A5A5A3", x"A2A29F9B", x"9A9B9B9B", x"9C99979A", x"9F9C9B9C", x"9B99999B", x"9D9B9895", x"94949799",
									 -- x"98989A9B", x"9C9FA1A3", x"A5A3A2A2", x"A4A7A8A9", x"A8ACB1B2", x"B1B1B3B5", x"B6B4B4B6", x"BABDBEBE",
									 -- x"C1BDBBBC", x"BDBDBEBF", x"C1C0BEBC", x"BCBAB8B6", x"B6B0AFB0", x"ADACADAC", x"A7A7A5A3", x"A3A4A4A3",
									 -- x"A2A3A3A2", x"A1A09F9F", x"A09E9C9B", x"9D9E9D9C", x"9F9E9D9E", x"A0A09E9C", x"9D9C9D9D", x"9E9D9A98",
									 -- x"9A98989A", x"9B9B9B9C", x"97999A9B", x"9A999898", x"9D9F9D9B", x"9D9C9A9C", x"9E9C9C9E", x"9E9D9D9E",
									 -- x"9D9D9D9B", x"9A9A9C9D", x"9C9D9EA0", x"A1A2A4A5", x"A8A7A6A5", x"A5A5A5A6", x"A6A5A5A7", x"ABADADAD",
									 -- x"A9AAAAAA", x"ABADB0B2", x"B3AEADAD", x"A8A7ABAC", x"A8AAABAA", x"ABADAFAF", x"ACADAEAF", x"B2B6BCC0",
									 -- x"C1C1C2C3", x"C4C6CBD1", x"D0D0CFCE", x"CCCACACA", x"CDCFCBC9", x"CAC4BFC3", x"C1C2C3C5", x"C6C6C9CC",
									 -- x"C6C6C6C7", x"C9C9C7C6", x"CBCDD0D2", x"D2D1D0CF", x"CFCFCFD0", x"D0CFCDCB", x"CDCDCCCA", x"C8C6C4C4",
									 -- x"C3C0BFC1", x"C0BBBABC", x"BDB7B3B5", x"B4B0AEAF", x"ACACABA9", x"A7A5A4A3", x"A3A5A7A7", x"A6A39F9C",
									 -- x"A0A3A29D", x"9B9C9C9A", x"9696938F", x"9194928D", x"8B8C8C8B", x"8A88827C", x"807C7979", x"7D818282",
									 -- x"7A858881", x"7C7B8089", x"9286817C", x"7F767776", x"74767571", x"6D69645E", x"615D5C5D", x"5B555457",
									 -- x"53595A54", x"53585B5A", x"62605E5A", x"5B63655E", x"5E5F5E61", x"5E5F6868", x"67686B6C", x"6B686666",
									 -- x"64605E61", x"625F5B59", x"5C5D5B59", x"585A5B5A", x"5B5B5C5E", x"5F5E5A58", x"59585654", x"53525252",
									 -- x"4B4E5153", x"52515152", x"57585958", x"58595A5B", x"5B5F6363", x"60606468", x"696B7074", x"787A7B7A",
									 -- x"7A7B7A79", x"787A7D7F", x"7E83878B", x"8E8D8E94", x"99979698", x"9C9E9C99", x"97999A99", x"999CA0A3",
									 -- x"A39F9B9A", x"98939191", x"8F92928B", x"8281807A", x"776F6B66", x"676A6362", x"5F5B5754", x"54545250",
									 -- x"504B4C4B", x"43434642", x"403D3A39", x"39373330", x"3131302F", x"2F302E2C", x"2B292828", x"29292724",
									 -- x"EAE9E8E7", x"E6E4E1E0", x"DAD5D1CE", x"CCC8C5C4", x"C3C3C1BF", x"BDBEC0C2", x"C4C5C5C5", x"C5C6C9CB",
									 -- x"CDCED0D3", x"D5D5D3D1", x"D2D3D1CD", x"CBCAC5BF", x"BFC0BDB9", x"B8B9B4AE", x"AFADACAD", x"AFAEABA7",
									 -- x"AAA7A5A6", x"A6A3A2A2", x"9F9E9D9C", x"9C9C9D9D", x"A1A2A09B", x"9B9D9C97", x"969B9B96", x"92939493",
									 -- x"9295989A", x"9B9C9E9F", x"9A9DA0A2", x"A4A8A9A7", x"A8ADAFB1", x"B4B3B2B4", x"B4B6B6B6", x"B8BCBEBE",
									 -- x"BCBDBDBD", x"BEC1C1C0", x"BFBFBFBF", x"BEBCBBBA", x"BAB3AEAF", x"AFACAAAB", x"AAA8A6A4", x"A3A3A3A2",
									 -- x"A4A3A2A0", x"9D9C9D9E", x"9F9E9C9C", x"9E9F9E9E", x"9F9D9EA1", x"A19E9FA3", x"A09FA09E", x"9C9FA19B",
									 -- x"999A9C9D", x"9D9B9A98", x"9C9C9B9A", x"999A9D9F", x"9E9D9B9B", x"9C9D9D9D", x"9F9E9E9F", x"A0A09F9E",
									 -- x"9F9FA0A0", x"9D9A9A9C", x"9C9B9C9F", x"A1A3A6A9", x"A6A7A6A5", x"A5A7A7A5", x"A6A6A6A7", x"A9AAABAB",
									 -- x"ACAAA9AA", x"ABACAFB2", x"B0AEACAB", x"A8A6A7AA", x"ABACABAA", x"ABADACA9", x"A9AEAFAC", x"ADB3B8B8",
									 -- x"B9BABDC0", x"C1C3C9CF", x"CFD1D0CD", x"CAC9C9C8", x"C8CCCDC8", x"C4C4C3C1", x"C4C3C2C3", x"C4C5C5C4",
									 -- x"C0C5C6C6", x"C7C6C5C8", x"CCCAC9CB", x"CED0D0CF", x"D0CFCFD0", x"CECBCACB", x"CAC9C8C8", x"C8C6C3C0",
									 -- x"C0C2C2BE", x"BBB9B8B6", x"B2B3B1AD", x"ACADADAB", x"AAA9A7A6", x"A5A4A3A2", x"A1A2A3A4", x"A3A09F9F",
									 -- x"9D9F9E9B", x"99999896", x"96909192", x"8D909490", x"8E8F8D88", x"8585837F", x"7C7D7D7E", x"8183827F",
									 -- x"7F7E7E80", x"7F7F8185", x"8283817D", x"79777572", x"75747372", x"6F6A6665", x"62605D5C", x"59585A5D",
									 -- x"5A5D645C", x"5D575E5F", x"65676765", x"65686969", x"66696665", x"68686769", x"6C6A6A6B", x"6E706F6D",
									 -- x"65655F63", x"5D605958", x"5F605F5C", x"5A5C5D5C", x"5A5B5F61", x"605D5C5F", x"5D5D5C5A", x"59585655",
									 -- x"50565955", x"50505356", x"59585859", x"595B6065", x"60656A6A", x"68676A6E", x"6D75787D", x"7F7E827F",
									 -- x"7D7D8084", x"84828387", x"86868F93", x"90929999", x"9D9E9FA0", x"A09F9F9F", x"A09EA2A2", x"9EA1A49D",
									 -- x"9FA0A19F", x"9C999797", x"918F8C8A", x"8885817E", x"75726D68", x"65635F5A", x"5B5C5A56", x"5351504F",
									 -- x"4C4B4A48", x"45434343", x"3F3B393A", x"39353230", x"2E2F2F2D", x"2B2B2B2A", x"2A292929", x"2A2A2826",
									 -- x"EBEAE8E6", x"E4E3E1DF", x"D8D4D0CE", x"CCC8C5C4", x"C1C2C1BF", x"BDBDBEBF", x"C2C3C4C3", x"C3C5C7C9",
									 -- x"CACBCCCF", x"D0D0CECC", x"D1D3D2D0", x"CFD0CCC6", x"C2C2C0BD", x"BCBDB9B2", x"B4B2AFAD", x"ADACACAB",
									 -- x"ABA7A5A6", x"A6A3A1A1", x"A2A2A09F", x"9F9FA0A0", x"A0A2A09C", x"9B9C9A95", x"959A9B96", x"93939290",
									 -- x"91939597", x"9898999A", x"9B9EA0A2", x"A4A7A8A7", x"A6ABADAF", x"B2B1B0B2", x"B3B5B6B6", x"B7BABBBA",
									 -- x"BDBEBDBC", x"BDC0C0BF", x"C0BFBFBF", x"BEBCBAB8", x"B7B1ADAF", x"AFADABAC", x"ABA9A6A5", x"A4A3A3A3",
									 -- x"A3A3A2A0", x"9F9E9FA0", x"9B9B9B9C", x"9D9E9D9C", x"9F9D9FA2", x"A29FA0A3", x"A09E9E9E", x"9C9FA19D",
									 -- x"9C9C9C9C", x"9C9C9C9B", x"9D9D9C9B", x"9A9A9C9E", x"9F9E9D9D", x"9C9D9E9E", x"A0A09FA0", x"A1A2A1A1",
									 -- x"A0A0A0A1", x"A09E9D9E", x"9D9C9D9E", x"9E9FA2A6", x"A5A6A5A4", x"A5A8A9A7", x"A8A6A4A5", x"A7A9A8A6",
									 -- x"ACAAA9AB", x"ABABADB0", x"AFAEADAC", x"A9A6A6A9", x"ABACACAC", x"ADAEADAB", x"AAADAEAD", x"AEB1B5B6",
									 -- x"B7B8BBBE", x"BFC1C6CB", x"CDCFCFCC", x"C9C8C8C7", x"C4C6C7C5", x"C3C3C2C2", x"C3C2C0BF", x"C0C2C3C3",
									 -- x"C1C4C4C3", x"C4C3C3C7", x"C4C7C9C9", x"C9C9CCCF", x"CDCDCDCC", x"CBC9C8C7", x"C8C6C5C5", x"C4C3C1BF",
									 -- x"BDBEBEBC", x"B9B8B6B4", x"B3B3B1AE", x"ACACABA9", x"A9A8A6A4", x"A4A4A4A3", x"A09FA0A1", x"A09E9EA0",
									 -- x"9C9D9C98", x"95959494", x"98929393", x"8E8F918C", x"8B8B8A87", x"8483807E", x"7D7D7C7C", x"7E81817F",
									 -- x"82818080", x"7E7D7E82", x"8182807C", x"79787674", x"72717070", x"6E6A6766", x"6362605F", x"5D5B5B5E",
									 -- x"5D5F6762", x"635E6568", x"666A6C6C", x"6C6D6C6B", x"6E706D6C", x"6E6D6C6D", x"6B6B6C6C", x"6B6B6B6B",
									 -- x"67676565", x"605F5C5C", x"5C5E5F5E", x"5E60605F", x"5B5C5F62", x"615F5F61", x"6161605E", x"5D5A5856",
									 -- x"56575758", x"5A5B5853", x"5F5C5A5A", x"5C5F6367", x"696C7071", x"706F7072", x"7579797D", x"7E7D8383",
									 -- x"82828486", x"86858688", x"8D8E9497", x"979BA0A2", x"A2A3A5A5", x"A3A3A5A7", x"AAA2A1A4", x"9F9A9B9F",
									 -- x"9D9E9E9D", x"9A979696", x"93908C88", x"85807C79", x"726F6A65", x"6464605C", x"57585652", x"50504E4C",
									 -- x"4A494745", x"44424140", x"3D3A3738", x"38353130", x"2F2F2E2B", x"2A2B2B2A", x"29292828", x"28292827",
									 -- x"ECEAE8E5", x"E3E1E0DE", x"D8D4D1D0", x"CDCAC7C6", x"C1C1C1C0", x"BEBDBDBD", x"C0C1C2C2", x"C2C2C4C6",
									 -- x"C8C9CBCD", x"CECECCCB", x"CCCFCFCF", x"D0D2CFCB", x"C6C7C6C3", x"C4C4C1BB", x"B9B7B4B1", x"AEADAEAF",
									 -- x"AEACA9A9", x"A8A6A4A3", x"A3A2A09F", x"9F9FA0A1", x"9FA1A09D", x"9C9B9792", x"93979996", x"9493918F",
									 -- x"90929495", x"96969696", x"9A9C9EA0", x"A2A5A7A7", x"A7ABADAE", x"B2B1B0B2", x"B1B3B4B5", x"B6B8B9B8",
									 -- x"BBBBBAB9", x"BBBEBFBE", x"C1C2C2C2", x"C1BFBCBA", x"B6B1AEAE", x"AFADACAC", x"AAA8A6A4", x"A3A3A2A2",
									 -- x"A1A1A1A0", x"9E9E9E9F", x"98999A9C", x"9D9D9B9A", x"9D9C9EA2", x"A2A0A0A3", x"A49F9FA1", x"9FA0A3A2",
									 -- x"A09F9D9C", x"9C9D9E9F", x"9F9F9F9E", x"9D9D9E9E", x"A0A0A09F", x"9D9D9FA0", x"A3A2A2A2", x"A3A3A3A3",
									 -- x"A09E9E9F", x"A09F9E9E", x"9D9D9D9D", x"9C9C9FA3", x"A4A4A4A4", x"A6A8A9A9", x"A8A5A3A4", x"A7A8A6A3",
									 -- x"AAA9AAAB", x"ACABACAD", x"AEADACAB", x"A8A5A5A7", x"AAACAEAD", x"ADAEAEAD", x"ADADAEAF", x"AFAFB2B5",
									 -- x"B4B5B8BB", x"BCBDC1C5", x"C9CCCCCA", x"C8C7C7C6", x"C5C4C2C2", x"C0BEBDBE", x"C0C0C0BF", x"BFBFC0C1",
									 -- x"C2C4C2C0", x"C2C2C2C7", x"C2C4C7C8", x"C8C8CACC", x"CACBC9C6", x"C6C7C6C2", x"C4C3C2C1", x"C0BFBEBE",
									 -- x"BBBBBAB8", x"B7B6B3B0", x"B0B0AFAC", x"AAA9A8A7", x"A7A5A3A2", x"A2A3A3A3", x"9F9E9D9D", x"9C9C9DA0",
									 -- x"9B9C9B97", x"93939494", x"938F9192", x"8F919390", x"8B898887", x"85817E7E", x"7E7E7C7A", x"7A7D7E7E",
									 -- x"81807F7E", x"7C7A7B7D", x"7E7E7D7A", x"77777573", x"71706F6F", x"6C686565", x"63626363", x"615E5F61",
									 -- x"60616767", x"6761676D", x"6F737678", x"78797876", x"74747372", x"72717070", x"6B6D6F6D", x"6A67686A",
									 -- x"68656461", x"63605F5B", x"585B5E5F", x"61626160", x"64646465", x"65626161", x"62626161", x"5F5D5A58",
									 -- x"5E5C5B5D", x"61635F59", x"625F5E61", x"6466696B", x"71747678", x"79787878", x"7F818085", x"8582898C",
									 -- x"8C8D8D8B", x"8B8B8A88", x"8F929496", x"9CA1A5A9", x"AAACADAB", x"A9A9ACB0", x"ADA9A6A6", x"A39B99A0",
									 -- x"A0A09F9D", x"9A989696", x"93908A85", x"807C7774", x"6F6C6763", x"6363605C", x"56555350", x"50504E4B",
									 -- x"48474443", x"42413F3D", x"3B383535", x"35333130", x"302F2C2A", x"2A2C2B29", x"28282827", x"27272829",
									 -- x"EBEAE8E6", x"E4E1DEDC", x"D9D5D2D1", x"CFCBC8C7", x"C4C3C1C1", x"BFBDBCBD", x"BFC0C1C1", x"C0C1C2C4",
									 -- x"C5C6C9CB", x"CCCDCCCC", x"C8CBCCCC", x"CED0CECB", x"C8C9C9C8", x"C8C9C7C3", x"BDBCB9B7", x"B5B3B2B1",
									 -- x"B2AFACAB", x"A9A7A5A4", x"A2A19F9E", x"9E9E9F9F", x"9E9F9F9C", x"9A999692", x"92949694", x"93939290",
									 -- x"91929395", x"95959595", x"98999A9C", x"9FA2A4A5", x"A8ABACAD", x"B1B1B0B2", x"B0B1B2B3", x"B5B7B8B9",
									 -- x"B6B7B6B6", x"B8BCBEBE", x"C0C1C2C2", x"C3C2BFBC", x"B7B3B0AF", x"AEACAAAA", x"A7A5A3A2", x"A2A2A1A1",
									 -- x"9F9F9E9D", x"9C9B9A9A", x"98999A9B", x"9C9B9A9A", x"9B9B9DA1", x"A2A0A0A2", x"A5A0A1A4", x"A3A2A3A4",
									 -- x"A1A09E9D", x"9D9EA0A1", x"A1A1A2A2", x"A2A1A1A1", x"A1A2A3A1", x"9F9FA1A3", x"A6A5A4A3", x"A3A3A4A4",
									 -- x"A19F9FA0", x"A09F9E9F", x"9C9D9E9F", x"9D9C9FA2", x"A2A2A3A4", x"A6A8A8A7", x"A6A5A5A6", x"A7A8A7A6",
									 -- x"A8A9AAAC", x"ADACABAB", x"ACACABA9", x"A6A5A5A7", x"A8ACAEAD", x"ACACACAC", x"ACAAABAF", x"AFACAEB2",
									 -- x"B2B3B5B8", x"BABABDC1", x"C5C8C9C8", x"C7C7C7C6", x"C8C4C1C1", x"C0BCBABC", x"BDC0C3C3", x"C1BFBEBD",
									 -- x"C0C2C0BE", x"C0BFC0C3", x"C3C3C3C5", x"C8C9C8C5", x"C6C8C5C1", x"C2C6C4BE", x"BFC0C0BF", x"BDBCBBBC",
									 -- x"BBBAB8B4", x"B3B2B0AC", x"ABABAAA9", x"A8A7A6A5", x"A3A2A1A0", x"A0A09F9F", x"A09D9B9A", x"99999C9F",
									 -- x"9C9D9C98", x"94949697", x"8E8C8D8E", x"8F929494", x"908B8888", x"86817E7F", x"7D7E7D7A", x"797A7B7A",
									 -- x"7C7C7C7A", x"78777779", x"797A7977", x"7575726F", x"6F6D6D6D", x"6B686767", x"63636465", x"64626264",
									 -- x"6665686A", x"69646972", x"797C7F82", x"83838383", x"78767777", x"74737372", x"6C6F716F", x"6B68696B",
									 -- x"6961605D", x"6764625B", x"5C5D5E60", x"62646463", x"6D6C6B6A", x"69686665", x"63616161", x"62605F5E",
									 -- x"60606060", x"61636464", x"6162666B", x"6F6F7072", x"76787C7D", x"7D7D7D7D", x"8587878F", x"8F898F93",
									 -- x"94969693", x"91918E89", x"8D929294", x"9FA5A7AD", x"AEAFAFAD", x"ABABAEB0", x"A6AFAEA8", x"A8A6A0A0",
									 -- x"A3A29F9D", x"9A979594", x"908C8681", x"7D797573", x"6D6A6662", x"62615D59", x"5554514F", x"4E4E4B47",
									 -- x"45454442", x"403F3D3C", x"39363333", x"3332312F", x"2F2E2B29", x"2A2C2B28", x"28282828", x"27252629",
									 -- x"EAE9E9E8", x"E6E2DEDB", x"DAD7D4D2", x"D0CCC9C7", x"C7C4C1C1", x"BFBCBCBD", x"BEBFC1C1", x"C0C0C1C2",
									 -- x"C2C3C5C7", x"C8C8C8C8", x"C8CACBCB", x"CCCDCBCA", x"C7C8C8C8", x"C9CBCAC8", x"C6C3BFBC", x"BBBAB7B4",
									 -- x"B4B2AEAA", x"A8A7A4A2", x"A3A2A1A0", x"A09FA0A0", x"9D9D9C9A", x"98979694", x"92929190", x"9091918F",
									 -- x"8F909192", x"93939493", x"9596979A", x"9C9FA2A4", x"A6A9A9AA", x"AEAEADAF", x"B0AFB0B1", x"B3B5B7B9",
									 -- x"B4B5B4B4", x"B6BABCBC", x"BCBEBEBF", x"C0C1BEBA", x"B8B4B1AF", x"ADABA9A8", x"A4A3A2A1", x"A1A1A1A0",
									 -- x"9D9D9C9B", x"99989797", x"98999998", x"98989898", x"999A9C9F", x"A0A0A0A0", x"A39FA1A5", x"A3A1A1A0",
									 -- x"A1A19F9E", x"9E9FA1A2", x"A1A2A3A4", x"A5A5A5A4", x"A3A4A5A3", x"A1A1A3A5", x"A5A5A4A4", x"A4A4A5A5",
									 -- x"A4A4A4A4", x"A19E9FA1", x"9D9EA0A1", x"A09E9FA1", x"A0A1A2A5", x"A6A6A5A4", x"A4A5A7A7", x"A6A6A7A8",
									 -- x"A7A8ABAC", x"ADADACAB", x"ABAAA8A5", x"A3A3A5A7", x"A6A9ABAA", x"A8A9A9A8", x"A8A5A6AB", x"ACA8A9AE",
									 -- x"B1B1B3B6", x"B8B8BBBE", x"C0C3C5C5", x"C5C6C6C6", x"C5C1BFC0", x"C1BEBEC1", x"BFC2C4C4", x"C2C0BEBE",
									 -- x"BDBFBDBC", x"BEBDBCBF", x"C1C0C0C2", x"C5C5C3C0", x"C3C5C3BF", x"C0C4C2BD", x"BBBCBDBD", x"BBB9B8B8",
									 -- x"BAB8B4B0", x"AFB0AEAC", x"A9A8A7A7", x"A6A4A3A3", x"A0A0A0A0", x"9F9E9C9A", x"9D9A9897", x"97979A9E",
									 -- x"9C9D9C98", x"94949596", x"8F8E8C8B", x"8D8F9092", x"948E8988", x"86817F7F", x"787B7C7B", x"7A7A7977",
									 -- x"77787877", x"75747576", x"76777776", x"74736F6B", x"6B696A6B", x"6C6B6B6C", x"67676869", x"67656668",
									 -- x"69686A6E", x"6C6C717B", x"7D808488", x"88868483", x"7E7A7B7C", x"76747574", x"6F70706E", x"6C6A6969",
									 -- x"68636460", x"68646560", x"63626264", x"66696B6C", x"6E6D6D6C", x"6D6D6C6A", x"68656365", x"66666667",
									 -- x"60626363", x"62636669", x"65696F74", x"7676787B", x"7C808283", x"807F8082", x"888A8A92", x"918B9195",
									 -- x"95999A98", x"9695928D", x"9097979A", x"A5ACADB1", x"AEADACAC", x"ADADADAD", x"A5AFAFA9", x"ABA9A3A1",
									 -- x"A09E9B99", x"97959290", x"8B87827D", x"79767371", x"6A686561", x"605F5A56", x"54524F4C", x"4B4A4642",
									 -- x"41424240", x"3D3B3A3A", x"38353231", x"3132302E", x"2C2C2A2A", x"2B2B2925", x"27272829", x"28252527",
									 -- x"EAEAEAEA", x"E9E5E0DD", x"DCD9D5D4", x"D2CECBC9", x"C9C5C2C1", x"C0BCBBBC", x"BEBFC1C1", x"C0C0C0C1",
									 -- x"C2C3C4C4", x"C4C3C4C4", x"C6C7C8C8", x"C8C8C7C7", x"C7C7C8C9", x"CBCDCDCD", x"D0CBC4C1", x"C0BFBCBA",
									 -- x"B9B6B2AD", x"AAA8A5A2", x"A2A2A2A1", x"A1A09F9F", x"9B9B9A98", x"96969696", x"93918F8D", x"8D8E8E8D",
									 -- x"8D8C8C8D", x"8E909090", x"95949699", x"9C9EA0A3", x"A4A7A6A7", x"ABACABAD", x"AFAEAEB0", x"B1B1B3B5",
									 -- x"B5B5B4B4", x"B5B8BAB9", x"BABCBCBB", x"BDBFBCB7", x"B5B3B0AE", x"ACAAA9A8", x"A4A3A2A2", x"A2A2A1A0",
									 -- x"9D9B9A99", x"98989796", x"97979695", x"94949597", x"99999B9D", x"9FA0A09F", x"A3A0A3A6", x"A4A3A3A0",
									 -- x"A2A1A1A1", x"A1A1A2A2", x"A2A2A3A5", x"A7A8A7A6", x"A6A7A6A5", x"A4A3A5A6", x"A3A3A4A4", x"A5A5A6A7",
									 -- x"A5A5A5A4", x"A19E9FA2", x"A0A0A1A2", x"A19F9E9F", x"A0A0A1A4", x"A6A5A3A3", x"A3A6A8A7", x"A4A3A4A6",
									 -- x"A6A8AAAB", x"ACADACAA", x"A9A9A7A3", x"A0A1A4A5", x"A5A7A7A6", x"A5A6A6A5", x"A7A4A5A9", x"AAA8A8AC",
									 -- x"AEAEB0B2", x"B4B5B8BB", x"BBBFC1C0", x"C0C2C3C3", x"C1C0BFBF", x"BFBEBFC1", x"C1C1C1C0", x"BFBEBFC0",
									 -- x"BCBEBDBC", x"BFBEBCBE", x"BEC0C3C3", x"C1BFBFC1", x"C0C1C0BE", x"BEC0BFBB", x"B8B9B9B9", x"B8B6B4B3",
									 -- x"B4B3B0AD", x"ACADADAB", x"A9A7A6A5", x"A3A1A0A0", x"9F9F9F9F", x"9F9C9997", x"97959494", x"9595989B",
									 -- x"9B9B9A96", x"93929290", x"8E8F8A88", x"8C8D8E92", x"948F8987", x"85817E7D", x"75777A7A", x"7A797774",
									 -- x"75767775", x"73737474", x"75767675", x"74736E6A", x"6C6B6A6B", x"6B6A6A6B", x"6D6D6D6E", x"6B69686A",
									 -- x"696A6A70", x"6E737983", x"7E81878B", x"89847E7C", x"80797B7C", x"73707472", x"71706E6C", x"6A686765",
									 -- x"64666865", x"64616566", x"68656467", x"6B6F7274", x"7071716F", x"6E6E6D6C", x"6F696668", x"6A69696B",
									 -- x"6766676A", x"6D6C6C6B", x"6F727679", x"797A7F85", x"86888987", x"84828486", x"8E908F92", x"908B9296",
									 -- x"94989B9B", x"99979593", x"989DA0A2", x"AAB0B2B3", x"AFAEADAE", x"B0B0AFAD", x"ACAAA7A7", x"A7A19EA1",
									 -- x"9C9A9796", x"9593908D", x"87837E79", x"75726F6D", x"6464625F", x"5C5B5855", x"52524F4C", x"49474440",
									 -- x"3D3E3E3D", x"3A383636", x"3634312F", x"2F302F2D", x"292A2A29", x"2A2A2724", x"27252629", x"28252426",
									 -- x"ECECECEC", x"EBE8E4E1", x"E0DCD9D7", x"D5D2D0CF", x"CCC7C4C5", x"C3BEBCBD", x"BDBFC1C1", x"C0BFBFBF",
									 -- x"C1C2C3C3", x"C2C1C2C3", x"C2C2C2C3", x"C3C3C4C5", x"C6C6C7C8", x"CBCDCFD1", x"D2CFCAC7", x"C5C4C1BF",
									 -- x"BEBBB6B0", x"ACAAA6A2", x"A1A1A2A2", x"A1A09E9D", x"9A9A9998", x"96949596", x"95928F8E", x"8F8F8E8D",
									 -- x"8D8C8A8B", x"8C8E8F90", x"94939598", x"9A9B9DA0", x"A2A4A2A3", x"A8A9A8AA", x"AAAAABAE", x"AFAEAEB0",
									 -- x"B3B3B3B2", x"B4B6B7B6", x"B7B8B8B8", x"BABEBBB6", x"B2B1AFAC", x"AAA9A7A6", x"A4A3A2A1", x"A1A09F9E",
									 -- x"9D9B9997", x"97969695", x"95959594", x"93939596", x"9A9A9A9C", x"9EA0A09F", x"A3A3A5A7", x"A5A6A6A1",
									 -- x"A3A3A2A2", x"A2A3A3A4", x"A4A4A5A7", x"A9ABAAA9", x"AAA9A8A6", x"A5A5A5A5", x"A3A4A5A6", x"A5A5A6A7",
									 -- x"A5A4A3A3", x"A19FA0A2", x"A19F9EA0", x"A09F9F9F", x"A1A0A0A3", x"A5A4A3A4", x"A3A6A7A7", x"A4A2A2A4",
									 -- x"A6A8A9A9", x"A9ABAAA9", x"A8A9A6A1", x"9FA0A1A2", x"A4A5A4A3", x"A3A5A5A4", x"A6A4A4A6", x"A7A7A7A9",
									 -- x"ABAAABAD", x"AFB1B4B7", x"B8BABCBB", x"BBBCBDBE", x"BEBFBFBC", x"BABABBBB", x"BEBDBBBA", x"BBBCBEBE",
									 -- x"BBBDBBBB", x"BEBDBBBD", x"BCBEC1C1", x"BEBDBEBF", x"BEBEBEBD", x"BCBBB9B8", x"B6B5B4B4", x"B4B2B0AE",
									 -- x"ADAEADAA", x"A9A9A9A8", x"A6A4A2A2", x"A09D9D9E", x"9D9D9D9C", x"9C999795", x"95939394", x"94939497",
									 -- x"98989795", x"9494918E", x"8C8E8988", x"8D8E8E93", x"908E8A86", x"84827E79", x"77777776", x"76767471",
									 -- x"71737472", x"71727372", x"74747372", x"72726E6A", x"6D6B6A6A", x"6A68686A", x"6E6E7071", x"6F6C6B6B",
									 -- x"6A6E6D73", x"6F777A81", x"7F818588", x"86807B79", x"7C737678", x"6D6C716F", x"716F6D6A", x"68676666",
									 -- x"63676768", x"6466676B", x"6A67686C", x"71747678", x"77797975", x"7271706E", x"736E6A6D", x"6E6D6D6E",
									 -- x"6F6D6E71", x"74747373", x"76787A7D", x"7E80858B", x"8C8B8A87", x"85858789", x"90959496", x"93909697",
									 -- x"989A9E9E", x"9B979799", x"9FA2A6A6", x"A8AEB1AE", x"B1B0B0AF", x"AFAFAEAD", x"ADA6A2A2", x"9F9D9E9D",
									 -- x"99969392", x"928F8B87", x"83807A76", x"726E6B69", x"6061605B", x"57565555", x"50504F4B", x"48464340",
									 -- x"3D3B3A39", x"39383532", x"3433302D", x"2E2F2D2A", x"28292928", x"27282624", x"26232326", x"27252427",
									 -- x"EEEDEEEE", x"EDEAE7E5", x"E3E0DCDB", x"D9D6D5D4", x"CEC9C7C9", x"C7C1BEBE", x"BDBFC1C1", x"C0BFBEBF",
									 -- x"BFC0C1C1", x"C0C0C1C2", x"C0BFC0C0", x"C1C2C4C6", x"C3C2C3C5", x"C7CACDD0", x"CECECECD", x"CBC8C5C3",
									 -- x"BFBDB7AF", x"ABA9A5A1", x"A1A2A3A3", x"A2A09F9D", x"9A999998", x"96949495", x"96939090", x"92929190",
									 -- x"908E8C8B", x"8D8F9191", x"93929397", x"99989A9C", x"9E9F9E9E", x"A3A4A3A5", x"A5A5A8AD", x"AEADACAD",
									 -- x"AFB0B0B0", x"B2B5B5B4", x"B1B3B3B3", x"B7BBBAB5", x"B1B0AEAB", x"A8A7A5A4", x"A4A3A1A0", x"A09E9D9C",
									 -- x"9E9C9896", x"95949392", x"94959595", x"94949597", x"9B9B9B9C", x"9EA0A09F", x"A2A3A5A4", x"A3A7A7A2",
									 -- x"A4A4A3A3", x"A3A4A5A5", x"A7A7A7AA", x"ACADADAC", x"ADABA9A7", x"A6A6A5A4", x"A5A6A7A7", x"A5A4A4A5",
									 -- x"A6A4A3A4", x"A4A3A3A4", x"A19D9B9D", x"9FA0A0A1", x"A2A0A0A2", x"A4A4A4A6", x"A4A5A6A6", x"A5A4A3A3",
									 -- x"A6A8A8A7", x"A7A9A9A7", x"A7A8A7A2", x"9E9F9F9F", x"A4A4A2A1", x"A3A6A6A4", x"A2A1A1A1", x"A2A3A3A4",
									 -- x"A8A6A7A9", x"ACAEB1B4", x"B5B8B9B7", x"B6B8B9B9", x"B9BDBDB9", x"B7B8B9B8", x"B8B7B7B8", x"BABBBBBA",
									 -- x"B8B9B7B6", x"BAB9B8BA", x"BBBAB9BA", x"BDBDBBB9", x"BDBCBCBD", x"BAB7B5B6", x"B5B3B0B0", x"B0AFADAB",
									 -- x"A9ACACA9", x"A7A5A5A4", x"A29F9E9E", x"9D9B9B9D", x"9A9A9999", x"98969493", x"96959596", x"94929293",
									 -- x"96979696", x"97989590", x"8C908B88", x"8E8E8C91", x"8E8E8B86", x"85847E77", x"7B797673", x"7373706D",
									 -- x"6C6F716F", x"6F717272", x"7373716F", x"6F706E6A", x"69676769", x"6A6A6C6E", x"6B6D7073", x"716E6C6D",
									 -- x"6F757376", x"7078787C", x"7F7F8081", x"7F7B797A", x"786E7275", x"6B6A7170", x"6F6E6C6A", x"68676868",
									 -- x"6767636A", x"69716E6F", x"6D6B6D72", x"7779797B", x"7A7D7F7C", x"78787776", x"77726F72", x"75737273",
									 -- x"71717273", x"7272757A", x"78797C80", x"8385898C", x"8C8A8785", x"8587898A", x"8C959799", x"97939795",
									 -- x"9E9FA1A2", x"9D97989D", x"A5A5A9A8", x"A5AAAFAA", x"B0B0AFAD", x"AAA9A9A9", x"A6A4A29C", x"99A0A297",
									 -- x"96938F8E", x"8C89837E", x"807C7873", x"706C6966", x"60615E58", x"53525354", x"4B4D4C49", x"46444240",
									 -- x"3F3B3738", x"3B3A3530", x"32322F2C", x"2D2E2C28", x"27292927", x"26262625", x"25202023", x"26242527",
									 -- x"F1F0EEED", x"EDEDEBE9", x"E6E2DEDA", x"D9D9D8D8", x"D2D0CAC6", x"C5C6C2BE", x"C1C2C3C3", x"C2C0BFBE",
									 -- x"C0BFBFBF", x"C0C0BEBD", x"BBBDBDBB", x"BCC0C1C1", x"BFBFC0C1", x"C4C7CACD", x"CBCDCDCB", x"CAC9C6C3",
									 -- x"C3BCB4B0", x"AEABA5A0", x"A5A3A2A0", x"A09F9E9D", x"99979695", x"93908F90", x"918F8F90", x"908F8F90",
									 -- x"8E8D8A8A", x"8D909190", x"92939395", x"979A9B9B", x"9A9B9C9F", x"A1A3A3A3", x"A5A7ABAD", x"AEADACAC",
									 -- x"B0AFAEAF", x"B1B2B1AF", x"AFB2B2AF", x"AFB3B5B4", x"B1AFADAC", x"AAA8A4A2", x"A4A4A2A0", x"9E9D9D9E",
									 -- x"9B979495", x"96949393", x"96929194", x"96969697", x"96999C9F", x"A0A0A1A2", x"A2A2A3A5", x"A5A4A4A6",
									 -- x"A5A4A4A4", x"A6A8A9A9", x"ABAAABAD", x"AEADADAE", x"ADADABAA", x"A8A8A8A9", x"ABA8A6A5", x"A6A7A6A4",
									 -- x"A3A3A4A5", x"A6A5A19E", x"9FA19F9E", x"A0A0A0A2", x"A4A2A1A3", x"A4A4A3A4", x"A5A3A3A4", x"A4A3A2A2",
									 -- x"9DA2A5A5", x"A4A6A5A3", x"A3A3A2A0", x"9F9FA2A4", x"A3A3A2A1", x"A1A2A09D", x"9FA0A1A1", x"A1A09F9F",
									 -- x"A4A5A7A9", x"ACAEB0B0", x"B4B5B6B6", x"B4B4B5B7", x"B6B4B3B3", x"B5B5B4B3", x"B5B3B1B2", x"B4B6B6B5",
									 -- x"B5B5B5B6", x"B7B7B7B6", x"B9BABCBB", x"B8B7B9BB", x"B9B5B5B8", x"B8B4B1B2", x"B0B4B3AD", x"A9ABABAA",
									 -- x"AAAAA9A8", x"A6A3A1A1", x"A09F9E9D", x"9D9C9A99", x"98999A99", x"95918E8C", x"90929492", x"8E8C8E90",
									 -- x"96979692", x"91929291", x"92908E8D", x"8E8F8E8E", x"8F8F8D87", x"817D7977", x"76777471", x"72706E70",
									 -- x"6D6F7170", x"6F706E6B", x"6C6D6D6D", x"6D6C6B6B", x"6C6A696B", x"69696E76", x"706F7172", x"7275746F",
									 -- x"6E747471", x"72737477", x"837D7776", x"7A7C7A77", x"72757671", x"6B696C70", x"65666A6E", x"6C67676B",
									 -- x"71706F70", x"73747270", x"7274777A", x"7F82807D", x"7A818786", x"817D7C7B", x"7D7A7777", x"78787673",
									 -- x"7873737A", x"7C79797D", x"80827F83", x"878A9394", x"8E87878B", x"8886898C", x"8E969992", x"969C9CA5",
									 -- x"A1A2A29F", x"9FA09F9C", x"9DA4A5A7", x"A7A6AAA7", x"AAA9A6A4", x"A5A7A6A4", x"9C9F9E9A", x"98999793",
									 -- x"918C8786", x"85807B77", x"75747371", x"6E6A6460", x"5D5B5754", x"5353504C", x"4B4A4744", x"4443403B",
									 -- x"403D3937", x"37373736", x"302F2E2E", x"2E2D2A28", x"282B2C29", x"24232424", x"23212124", x"27262524",
									 -- x"F1F1F1F1", x"F0EFEDEB", x"E7E5E1DF", x"DDDCDBD9", x"D7D4CEC9", x"C7C7C3BF", x"C0C1C2C2", x"C1BFBEBD",
									 -- x"BEBDBDBD", x"BEBEBCBB", x"B9BBBCBB", x"BCBFBFBE", x"BEBEBEBF", x"C1C5C9CC", x"CCCDCCCA", x"C9C7C4C1",
									 -- x"C2BDB8B5", x"B3B0ABA6", x"A3A2A1A0", x"9F9E9B9A", x"96949292", x"918E8E8F", x"8E8D8D8E", x"8E8E8F90",
									 -- x"8C8A8888", x"8B8E9090", x"94949495", x"97999A9A", x"9A9A9B9D", x"9FA1A1A1", x"A2A3A4A5", x"A6A7A9AA",
									 -- x"ACABAAAC", x"AEAFAEAD", x"AEAFAEAC", x"AEB2B2AF", x"ACAAA8A7", x"A6A5A3A1", x"A3A3A2A1", x"A09F9F9E",
									 -- x"9B989696", x"96949495", x"95939295", x"9797989A", x"989A9DA0", x"A1A1A1A2", x"A0A1A3A5", x"A6A4A4A5",
									 -- x"A8A8A8A8", x"A8A8A9A9", x"AAA9ABAF", x"B0B0B0B1", x"B0ADA9A9", x"ABABA8A5", x"ABA9A7A7", x"A7A8A7A6",
									 -- x"A3A3A3A5", x"A6A5A2A0", x"A2A4A19E", x"9F9FA0A4", x"A4A3A4A5", x"A4A2A2A3", x"A1A0A0A1", x"A2A09E9E",
									 -- x"A1A2A2A1", x"A0A2A3A3", x"A5A3A09D", x"9B9B9EA0", x"A09F9E9D", x"9D9E9D9B", x"999B9C9D", x"9D9D9D9D",
									 -- x"9F9E9FA3", x"A8ABADAC", x"ACAEAFB1", x"B1B2B3B4", x"B1AFADAE", x"B0B0B0AF", x"B2B1B0B0", x"B2B3B4B4",
									 -- x"B3B3B4B6", x"B7B7B6B4", x"B7B7B7B8", x"B8B7B6B6", x"B3B0B0B4", x"B4B0AFB1", x"ADAEAEAB", x"AAAAAAA9",
									 -- x"A8A6A4A2", x"A1A1A1A2", x"A1A09F9D", x"9B989593", x"97979695", x"93918F8D", x"8D8F9090", x"8F909193",
									 -- x"92939290", x"8F929494", x"9090908E", x"8C8B8C8E", x"8B8C8B87", x"83817F7D", x"7A7A7571", x"716E6B6D",
									 -- x"6B6E6F6E", x"6F706F6D", x"6D6C6B6B", x"6A6A6A6A", x"6D6A686B", x"6C6C7177", x"77737577", x"76767672",
									 -- x"72777774", x"7678787B", x"7F7B7777", x"797A7876", x"7674716F", x"6E6E6D6D", x"6A6A6D70", x"6F6C6C70",
									 -- x"7174787A", x"7B7A7877", x"747B8284", x"85868889", x"7F858989", x"87878889", x"85837F7D", x"7D7B7977",
									 -- x"7877787B", x"7E808080", x"8789868A", x"8D8E9594", x"918B8A8A", x"8584898D", x"91939796", x"9DA5A3A5",
									 -- x"A2A2A19D", x"9D9FA1A1", x"A1A6A3A3", x"A3A3A9A7", x"A7A7A6A5", x"A4A5A4A2", x"9C9D9B98", x"98999690",
									 -- x"8F898380", x"7E7A7573", x"716E6B67", x"6563605E", x"57575551", x"4F4F504F", x"4E4A4440", x"3F3F3E3B",
									 -- x"3C393534", x"34353434", x"312F2D2D", x"2D2C2A28", x"28292926", x"24242423", x"22201F22", x"24242323",
									 -- x"F2F3F4F3", x"F1EFEDEC", x"E9E8E6E4", x"E3E1DEDC", x"DBD8D2CD", x"CBC9C6C2", x"C0C1C1C1", x"C0BEBDBC",
									 -- x"BCBCBBBB", x"BCBCBBBA", x"B6B9BABB", x"BCBDBCBB", x"BFBFBFBF", x"C1C5C9CD", x"CACBCBC8", x"C6C5C2C0",
									 -- x"BEBCB9B8", x"B5B2ACA8", x"A2A1A0A0", x"9F9E9B99", x"9391908F", x"8E8D8E8F", x"8D8B8A8B", x"8C8C8D8F",
									 -- x"8C8A8889", x"8B8E9091", x"93939394", x"9697999A", x"9999999A", x"9C9D9E9E", x"9FA0A0A1", x"A2A4A6A8",
									 -- x"A9A8A9AA", x"ACADACAA", x"AAAAAAA9", x"ADB1B0AC", x"AAA8A5A4", x"A3A3A2A1", x"9F9E9E9E", x"9F9E9D9B",
									 -- x"9B9A9998", x"96959597", x"95949596", x"9697989A", x"9A9C9FA1", x"A2A2A2A2", x"A1A1A4A7", x"A7A5A5A6",
									 -- x"AAABACAC", x"ABAAABAC", x"ACACADB1", x"B3B3B3B3", x"B1AFADAC", x"ADACA9A6", x"A9A9A8A7", x"A7A7A7A7",
									 -- x"A3A2A2A4", x"A5A6A4A3", x"A3A5A29E", x"9D9D9FA6", x"A2A3A4A5", x"A29F9FA1", x"9F9E9E9F", x"A09E9D9D",
									 -- x"A19F9E9F", x"A0A0A1A3", x"A4A3A09D", x"9B9B9B9D", x"9C9C9A99", x"9A9B9B99", x"97989A9B", x"9B9B9C9D",
									 -- x"9C9A9A9D", x"A3A8A8A7", x"A8A9AAAD", x"AFB0B1B0", x"AEACAAAA", x"AAACABAB", x"AAABACAC", x"ADAEB0B1",
									 -- x"AFAFB0B1", x"B2B3B3B3", x"B3B2B2B4", x"B6B5B3B0", x"B3B1B0B1", x"AFABAAAC", x"AAA7A6A8", x"AAA9A7A7",
									 -- x"A7A4A09F", x"9FA1A1A0", x"9C9C9C9C", x"9B999694", x"96949291", x"9291908F", x"8B8C8C8D", x"8E8F9091",
									 -- x"8C8D8D8C", x"8C8E9090", x"8F91928F", x"8A888A8D", x"898A8984", x"807E7B79", x"7777736F", x"706F6D70",
									 -- x"6B6D6F6F", x"6F6F6F6E", x"6E6D6B6A", x"6A6C6D6E", x"706C6B6F", x"7274777B", x"7C767679", x"78767776",
									 -- x"787A7674", x"77797A7D", x"7C7B7A79", x"79787776", x"77747170", x"71716F6D", x"6E6D6E71", x"72707174",
									 -- x"777B8184", x"83828182", x"8486888B", x"8D8F8D89", x"90929390", x"8D8B8A88", x"8B898684", x"827F7D7C",
									 -- x"7B7E7F80", x"84898A87", x"8C908E92", x"93919593", x"938F8E8A", x"84868D8F", x"8F8B9195", x"9DA8A49F",
									 -- x"A5A5A3A0", x"9FA1A2A3", x"A5A9A5A5", x"A3A3A8A7", x"A2A4A4A2", x"A1A1A09E", x"9B9B9895", x"9595918A",
									 -- x"88837E7C", x"7B777371", x"6E6B6763", x"605E5D5C", x"5557554F", x"4B4A4B4C", x"4F4B4540", x"3E3E3D3A",
									 -- x"37353231", x"3131302F", x"302E2C2B", x"2B2A2927", x"26272624", x"23242422", x"24211F21", x"22222324",
									 -- x"F4F5F5F3", x"F0EDEBEB", x"EBEAE9E8", x"E8E5E2DF", x"DDDAD5D1", x"CDCBC8C6", x"C2C2C1C1", x"C0BEBCBB",
									 -- x"BBBBBBBB", x"BBBBBBBA", x"B6B8B9BA", x"BBBBBAB9", x"BEBFBFC0", x"C2C5C9CB", x"C8C9C9C7", x"C4C3C1BF",
									 -- x"BBBBBAB9", x"B6B1ABA7", x"A4A2A09F", x"9F9E9C9A", x"93918F8F", x"8E8D8E90", x"8C8A898A", x"8989898B",
									 -- x"8D8A8888", x"898B8C8E", x"908F9092", x"94959799", x"98979797", x"98999A9A", x"9A9B9EA0", x"A1A2A2A3",
									 -- x"A5A5A6A8", x"A9A9A8A7", x"A5A7A7A8", x"ABAFAEAB", x"ABA8A4A2", x"A1A1A09F", x"9D9B9A9A", x"9C9D9B99",
									 -- x"9A9B9B9A", x"97959697", x"95969796", x"95959699", x"9C9EA0A2", x"A3A3A3A2", x"A3A3A5A7", x"A8A7A7A9",
									 -- x"AAADB0B1", x"B0AFAFB1", x"B1B1B2B4", x"B5B4B3B2", x"B0B2B4B2", x"AEAAAAAB", x"A8A8A8A7", x"A6A5A4A5",
									 -- x"A3A2A2A3", x"A4A5A6A5", x"A1A3A09C", x"9B9A9DA5", x"A1A1A2A3", x"A29F9E9F", x"9E9B9A9B", x"9C9B9B9C",
									 -- x"9B98999E", x"A09E9D9E", x"9D9E9E9E", x"9D9B9998", x"99989796", x"97989795", x"95969898", x"9899999A",
									 -- x"9998989A", x"9EA1A1A0", x"A5A5A7A9", x"ACADACAB", x"ACAAA8A5", x"A5A6A6A5", x"A2A4A7A7", x"A7A7AAAC",
									 -- x"ACABA9AA", x"ABADAFB0", x"B0AFAEB0", x"B1B1AFAD", x"B1AFAFAF", x"ABA8A7A9", x"A8A2A0A5", x"A9A6A3A4",
									 -- x"A6A4A1A0", x"A1A29F9B", x"99999B9C", x"9C9B9896", x"95929090", x"9191908F", x"8C8C8C8B", x"8A898A8B",
									 -- x"8C8C8C8C", x"8B8B8C8C", x"9192908C", x"8785878A", x"8888847F", x"7B797775", x"7475716E", x"706F6F72",
									 -- x"6C6E7070", x"6F6E6D6D", x"6F6E6E6E", x"6F717375", x"74737477", x"7B7C7E80", x"817A797D", x"7A78797A",
									 -- x"7E7D7774", x"777A7B7E", x"7D7D7D7C", x"7A797979", x"75767674", x"72717172", x"71707174", x"76767679",
									 -- x"7E818589", x"89898A8C", x"90909090", x"9293918D", x"95989A9A", x"9997938F", x"8F8E8C89", x"87858484",
									 -- x"81828588", x"8D919291", x"92969598", x"98959692", x"918E8D89", x"868A8F8F", x"8D879095", x"9BA6A49D",
									 -- x"A6A6A6A5", x"A5A3A09E", x"A4A8A7A9", x"A8A3A4A0", x"9C9FA09D", x"9B9A9A99", x"9A999590", x"8F8E8984",
									 -- x"827E7C7B", x"79746E6A", x"69686664", x"605D5A58", x"5657554F", x"4A494949", x"49484541", x"403E3B37",
									 -- x"36343231", x"302E2C2A", x"2E2D2B2A", x"2A292725", x"25252523", x"22232322", x"25211F20", x"20212224",
									 -- x"F6F6F5F2", x"EFEDECED", x"EEECEBEA", x"EAE8E4E2", x"DFDCD8D4", x"D0CCC9C8", x"C4C3C2C1", x"C1BFBDBB",
									 -- x"BBBBBBBA", x"BABABABA", x"B8B8B9BA", x"BBBABABB", x"BCBDBFC1", x"C2C4C6C7", x"C7C9C9C6", x"C2C1BFBD",
									 -- x"BBBBBCBB", x"B8B3AEAA", x"A7A4A09E", x"9D9D9A98", x"94918F8F", x"8E8C8D8F", x"8B898889", x"88878889",
									 -- x"8A868484", x"8586888B", x"8F8E8F91", x"92929599", x"96959393", x"94959696", x"95979A9C", x"9D9D9E9E",
									 -- x"9E9FA0A2", x"A4A4A4A3", x"A4A6A8A8", x"A9AAABAA", x"A8A6A3A0", x"9F9F9D9C", x"9D9B9999", x"9A9B9A99",
									 -- x"979A9C9B", x"98969697", x"95979997", x"9596989A", x"9D9EA0A2", x"A4A4A3A2", x"A5A5A5A7", x"A8A8AAAC",
									 -- x"ACB0B3B5", x"B4B3B4B5", x"B7B6B6B6", x"B7B6B4B1", x"B2B4B5B3", x"AFABABAD", x"A9AAAAA8", x"A6A4A3A3",
									 -- x"A3A3A2A2", x"A3A4A5A6", x"A0A2A09D", x"9C999BA3", x"A3A0A0A2", x"A3A29F9E", x"9C989696", x"96969799",
									 -- x"9896979B", x"9D9A9899", x"98989999", x"99979593", x"95959493", x"94949390", x"92929394", x"94949596",
									 -- x"92939597", x"97989999", x"A0A0A1A3", x"A6A7A6A4", x"A5A5A39F", x"9FA0A19F", x"9FA1A4A4", x"A2A2A3A5",
									 -- x"A6A5A5A6", x"A8AAABAB", x"ABACACAC", x"ACABACAC", x"A8A9A9A9", x"A7A6A6A8", x"A7A09DA2", x"A5A29FA0",
									 -- x"A6A4A1A0", x"A2A3A09A", x"9C9C9C9C", x"9C999694", x"9492908F", x"90908E8C", x"8C8D8E8B", x"87858689",
									 -- x"8F8E8C8B", x"8B8C8E91", x"93918E89", x"85848586", x"8584817D", x"7B7B7B79", x"7777736F", x"6F6E6C6E",
									 -- x"6A6D7072", x"706E6D6D", x"6F707173", x"75767778", x"797A7D81", x"82828385", x"8A828184", x"817D7F80",
									 -- x"83827D7C", x"7F807F81", x"80807F7D", x"7B7A7A7B", x"77777675", x"74737474", x"7676777A", x"7C7D7D7E",
									 -- x"8283878D", x"91929293", x"90989D99", x"9392979C", x"9C9EA1A2", x"A4A39F9A", x"97969390", x"8D8B8A8A",
									 -- x"88868990", x"95959699", x"999D9B9F", x"9E999995", x"8E8B8B8A", x"8A8E8F8A", x"8F8B969A", x"9DA6A8A5",
									 -- x"A7A5A4A5", x"A6A39E99", x"9FA3A4A8", x"A69F9E99", x"999B9B98", x"95959594", x"9695928D", x"89878482",
									 -- x"7F7B7877", x"736D6763", x"63636260", x"5D5A5655", x"5252504D", x"4C4B4A47", x"4142413E", x"3D3C3835",
									 -- x"35343332", x"302E2C2A", x"2B2A2929", x"29282523", x"23262623", x"20212223", x"24211E1E", x"1E1E1F22",
									 -- x"F7F6F5F3", x"F1F0F1F1", x"EFEEEDED", x"ECEAE7E4", x"E1DFDCD8", x"D2CCC9C9", x"C7C5C3C2", x"C2C0BEBC",
									 -- x"BABABABA", x"B9B9BABA", x"BCBBBABB", x"BCBBBBBD", x"BDBFC1C2", x"C3C4C5C6", x"C8CAC9C5", x"C1BFBDBC",
									 -- x"BABABAB9", x"B8B4B0AD", x"AAA6A09D", x"9B9A9794", x"93918F8E", x"8D8B8C8D", x"89888889", x"8988888A",
									 -- x"87848283", x"8484878B", x"8F8E8E90", x"908F9297", x"93929190", x"91929292", x"95959697", x"98999B9D",
									 -- x"98999B9E", x"A0A1A2A2", x"A4A5A6A6", x"A5A5A6A7", x"A5A3A1A0", x"A09F9D9B", x"9B999796", x"97979797",
									 -- x"95989A99", x"98979796", x"96989A99", x"989A9C9D", x"9E9FA1A3", x"A5A5A4A3", x"A6A5A5A7", x"A8A9ADB0",
									 -- x"B2B4B7B9", x"B9B8B7B8", x"BAB9B8B8", x"B9BAB8B5", x"B7B4B1B0", x"B1B0ADAB", x"ADACACAB", x"AAA7A5A4",
									 -- x"A5A4A3A2", x"A2A3A4A5", x"A2A2A09F", x"9E9A9AA1", x"A6A2A0A2", x"A5A3A09E", x"9C989595", x"95959698",
									 -- x"9D9A9999", x"9998999A", x"99979593", x"93939392", x"94949392", x"9293918E", x"8F8F9091", x"91929393",
									 -- x"8D909293", x"93939596", x"999A9B9E", x"A0A1A1A1", x"9EA09F9B", x"9B9E9F9E", x"9EA0A2A2", x"A09E9E9F",
									 -- x"9FA1A3A6", x"A8A7A5A4", x"A6A8A9A8", x"A6A5A7AA", x"A6A7A7A6", x"A5A4A3A3", x"A49F9C9F", x"A09D9D9F",
									 -- x"A4A39F9D", x"A0A3A29E", x"9E9D9D9C", x"9B999795", x"94939191", x"908F8C8A", x"8C8E8F8C", x"88878A8D",
									 -- x"8F8C8887", x"888B9196", x"96938E8B", x"89888786", x"83827F7B", x"7A7B7A78", x"77787572", x"726F6C6E",
									 -- x"696C7073", x"73717072", x"72737679", x"7B7B7A79", x"7F818587", x"87878889", x"928C8B8B", x"87858788",
									 -- x"88898788", x"8B898587", x"8583817F", x"7E7E7D7C", x"7C797676", x"797B7976", x"7A7B7D7F", x"80818384",
									 -- x"85868B96", x"9C9C9998", x"979D9F9C", x"98989B9F", x"A3A5A6A7", x"A9AAA7A4", x"A09D9894", x"918F8D8C",
									 -- x"908C8F98", x"9C9A9B9F", x"9EA19FA2", x"A19B9B96", x"928D8D8F", x"9091908A", x"8E8D979A", x"9EA6A7AA",
									 -- x"AAA6A2A3", x"A3A19E9C", x"9DA09EA2", x"A19B9B97", x"96979693", x"9191908F", x"8F8E8C89", x"86838180",
									 -- x"7B777371", x"6E6B6867", x"60605E5B", x"58565656", x"51504D4A", x"4A494540", x"403F3D3A", x"393A3937",
									 -- x"33333231", x"302E2D2C", x"29282727", x"28272422", x"22252623", x"1F202224", x"2522201F", x"1F1E1F21",
									 -- x"F7F6F5F4", x"F4F4F3F3", x"F1F0F0F0", x"EFEDE9E6", x"E3E1DFDC", x"D6CFCBCB", x"C9C7C4C3", x"C2C1BEBC",
									 -- x"BABBBBBA", x"BABABBBC", x"BEBDBDBE", x"BEBDBDBF", x"C0C1C3C4", x"C4C5C5C6", x"C7C9C9C5", x"C1BFBEBD",
									 -- x"BCBAB8B7", x"B6B3AFAC", x"ABA7A19D", x"9C9A9693", x"92908F8E", x"8D8B8B8D", x"8988888A", x"8A898889",
									 -- x"88848283", x"8483878C", x"8D8B8B8E", x"8D8C8F94", x"908F8E8E", x"8F8F8F8F", x"91929394", x"94959798",
									 -- x"9597999B", x"9C9E9FA0", x"A2A1A1A1", x"A1A2A2A3", x"A1A09F9F", x"9F9E9B99", x"96969594", x"94949494",
									 -- x"94979896", x"96979796", x"97999A99", x"999C9E9E", x"A0A0A2A4", x"A6A7A6A4", x"A5A5A6A9", x"ABAEB1B5",
									 -- x"B7B8BBBC", x"BDBCBBBA", x"BDBCBABA", x"BCBEBDBA", x"BAB6B1B0", x"B2B2B0AD", x"AFAEAEAD", x"ADABA8A5",
									 -- x"A6A5A4A2", x"A1A1A2A2", x"A2A19F9F", x"9F9C9CA3", x"A7A4A2A3", x"A3A19E9C", x"9C999796", x"96959597",
									 -- x"9C9B9995", x"94959798", x"98969391", x"91919191", x"91918F8D", x"8E908F8D", x"8D8E8E8E", x"8E8E8F8F",
									 -- x"8C8D8D8E", x"8E909293", x"92949698", x"999A9B9C", x"999B9B98", x"989C9D9B", x"9A9C9E9E", x"9D9C9C9C",
									 -- x"9B9D9FA2", x"A3A3A19F", x"A0A3A5A4", x"A2A1A2A4", x"A7A6A5A4", x"A3A19E9C", x"A09D9B9B", x"9A9A9CA0",
									 -- x"A1A2A09E", x"A0A5A4A0", x"A1A09E9E", x"9D9D9C9B", x"98979694", x"92908E8D", x"8E8F8F8D", x"8B8A8D8F",
									 -- x"8B888686", x"87898D92", x"92908D8C", x"8B898785", x"81807E7B", x"7A797673", x"75777675", x"76737071",
									 -- x"6D6F7377", x"7776787B", x"777A7D81", x"83828180", x"8788898A", x"8C8D8E8D", x"96939393", x"90919493",
									 -- x"95959392", x"94918E91", x"8F8B8786", x"87878481", x"827F7C7C", x"7F80807E", x"7F818383", x"8385888A",
									 -- x"8F8F949E", x"A4A29E9D", x"9F9F9E9E", x"A0A2A19E", x"A0A4A8AC", x"B0B2B1AF", x"A4A09A96", x"95949392",
									 -- x"9897999F", x"A3A3A3A4", x"A3A5A2A4", x"A29D9D99", x"97908F93", x"9392918F", x"8E8E9396", x"9FA5A3A7",
									 -- x"A9A5A2A0", x"9E9B9A9C", x"9A9B979B", x"9A969896", x"9292918F", x"8E8D8B88", x"87868585", x"83807C79",
									 -- x"76726F6E", x"6C6A6868", x"605F5C59", x"55535354", x"524F4B47", x"45443F3A", x"403F3C38", x"37383837",
									 -- x"31313130", x"2F2D2C2C", x"29272525", x"25252524", x"21232321", x"1F212324", x"26242322", x"211F2021",
									 -- x"F7F6F5F5", x"F5F4F2F1", x"F2F2F2F2", x"F2EFEBE7", x"E3E2E1DF", x"D9D1CECF", x"C9C7C4C3", x"C3C1BFBC",
									 -- x"BCBDBDBC", x"BBBBBCBE", x"C0BEBEC0", x"C0BEBEC0", x"C1C1C2C2", x"C2C3C4C5", x"C5C7C8C4", x"C1C0C0C0",
									 -- x"C0BDB9B6", x"B5B3AFAC", x"AAA6A19F", x"9E9C9894", x"92908F8F", x"8F8D8C8D", x"8A898A8B", x"8B888788",
									 -- x"88848182", x"82808489", x"8887888A", x"8A898D93", x"8F8E8D8D", x"8E8E8E8E", x"8A8D9092", x"92919090",
									 -- x"93949697", x"98999A9B", x"9F9D9A9C", x"9EA0A1A1", x"9D9C9C9C", x"9C9A9694", x"95969696", x"95959595",
									 -- x"94969694", x"94969897", x"989A9A99", x"999C9D9D", x"A1A1A2A5", x"A7A8A7A5", x"A5A5A8AC", x"AFB2B5B9",
									 -- x"BABABCBE", x"C0C0BFBD", x"BFBEBCBB", x"BDC1C0BC", x"BAB9B6B3", x"B2B1B3B4", x"B0AEADAE", x"AEADA9A6",
									 -- x"A7A6A4A2", x"A0A0A0A1", x"A09F9C9D", x"A09E9FA6", x"A7A5A3A2", x"A09C9A9A", x"9A989696", x"95949394",
									 -- x"93969590", x"8E919392", x"9391908F", x"90908F8E", x"8C8B8886", x"878A8B8A", x"8B8B8B8A", x"89888989",
									 -- x"8C8A8887", x"898B8D8E", x"8D8F9191", x"92929496", x"94989895", x"94989896", x"9496999B", x"9C9C9B9B",
									 -- x"9B9A9B9C", x"9D9E9E9D", x"9C9FA1A2", x"A09F9FA0", x"A1A1A0A0", x"A09F9C99", x"9C9C9A98", x"96989CA1",
									 -- x"9FA2A3A2", x"A4A7A49E", x"A6A5A2A0", x"9F9F9E9D", x"9C9B9A97", x"94929292", x"92918F8D", x"8C8C8C8D",
									 -- x"8988898B", x"8B88888A", x"89898989", x"88858381", x"7E7E7E7C", x"7B7A7672", x"76797877", x"78757172",
									 -- x"7274777B", x"7B7A7D82", x"7C7F8387", x"8A8A8988", x"8E8C8A8B", x"8F929291", x"98989A99", x"989CA09F",
									 -- x"A6A39D9A", x"9A97979C", x"97938E8E", x"908F8B86", x"84858684", x"82828588", x"85878988", x"87898E91",
									 -- x"9A989BA3", x"A7A4A2A2", x"9CA1A4A5", x"A6A7A9A9", x"A9AEB3B5", x"B6B4AFAA", x"A6A19B99", x"9A9B9B9A",
									 -- x"9EA0A2A5", x"A8ACABA8", x"A8AAA6A7", x"A59FA09C", x"968E8E93", x"918F9091", x"94939496", x"A3A8A1A5",
									 -- x"A4A2A09D", x"97929295", x"95959195", x"95919392", x"8E8E8D8C", x"8B8A8783", x"82807F81", x"817D7671",
									 -- x"74716E6D", x"6A65615F", x"5E5D5B57", x"534F4E4D", x"4F4D4945", x"4342403C", x"3D3D3A37", x"35353533",
									 -- x"3030302F", x"2D2B2A29", x"29262422", x"23242525", x"2122211F", x"20222423", x"24232222", x"201E1E20",
									 -- x"F4F5F6F6", x"F5F4F3F3", x"F6F4F2F0", x"EFEEECEB", x"E3E2DFDB", x"D8D6D3CF", x"CBC8C7C7", x"C5C1BEBE",
									 -- x"C2C0BEBD", x"BDBEBEBE", x"C1C1C0C0", x"C1C1C0C0", x"C2C2C2C1", x"C0C0C1C1", x"C3C4C5C4", x"C2C1C0C1",
									 -- x"C1BEBAB7", x"B5B2ADA9", x"A7A29E9D", x"9F9F9A95", x"92908F8F", x"8F8D8D8F", x"8B8B8C8C", x"8B8A8887",
									 -- x"86868584", x"84848485", x"85888987", x"888B8E8F", x"8C8D8D8C", x"8B8B8C8D", x"8D8B8B8C", x"8C8D8F92",
									 -- x"938F8E93", x"97969698", x"999E9E98", x"979B9C99", x"9D9B9998", x"99999795", x"94939293", x"94959492",
									 -- x"90949899", x"99989694", x"9A979698", x"9C9F9F9D", x"9FA0A4A8", x"A9A8A9AB", x"ABABABAE", x"B2B8BEC1",
									 -- x"BFBEBFC2", x"C2C1C0C1", x"C1C3C2BE", x"BCBFC1C2", x"BBBCB7B2", x"B6B8B4B0", x"B0B0AFAE", x"AEACA9A6",
									 -- x"A6A7A7A5", x"A5A6A4A1", x"A0A0A0A0", x"9F9D9EA1", x"A5A7A7A4", x"9F9D9B99", x"98989694", x"9494928F",
									 -- x"90909090", x"90919090", x"90908F8F", x"8E8C8A89", x"898B8A86", x"83838382", x"87898885", x"84868683",
									 -- x"88858486", x"8686888B", x"878C878C", x"8E8C9490", x"90929494", x"93919091", x"96949696", x"93959A9A",
									 -- x"96989A9B", x"9B9B9B9C", x"999B9D9E", x"9D9D9D9E", x"9E9B9B9E", x"9E9B9A9C", x"989CA09F", x"9C9A9DA0",
									 -- x"A3A4A7AA", x"A8A5A5A8", x"A6A4A2A3", x"A5A5A29F", x"A4A29E9B", x"99989696", x"96938F8E", x"8D8D8A88",
									 -- x"868A8687", x"8B8E9089", x"918B8288", x"8882857C", x"7D7D7C7B", x"7A787879", x"77777775", x"74747678",
									 -- x"73777B7E", x"7F828689", x"85848C93", x"90909392", x"94959596", x"989B9C9C", x"9A9EA4A6", x"A4A0A3A9",
									 -- x"AFAEADA9", x"A29D9EA3", x"A0A3A29A", x"9594918C", x"878E8C88", x"8D8D8A8D", x"8E93918E", x"9094979C",
									 -- x"9B9D9EA0", x"A5A9A59D", x"A3A4A6A8", x"AAAAA8A6", x"A8B3B2B8", x"C2C2BBB2", x"ACA1A0A5", x"A4A7A8A1",
									 -- x"A4A6A7A6", x"A6A9ABAC", x"AEB0AFAB", x"A8A6A099", x"99979491", x"8F8F9091", x"9093979D", x"A4A8A7A4",
									 -- x"A19A999A", x"98969593", x"92929190", x"93959694", x"8F8C8887", x"88898784", x"82807D7B", x"79787674",
									 -- x"706D6A68", x"6765605D", x"5B575556", x"55504D4B", x"4F4C4947", x"443F3C3D", x"3B3A3836", x"35353330",
									 -- x"332F2E30", x"2F2B2829", x"2D2A2725", x"24242322", x"22211F1F", x"1F212223", x"21201F1D", x"1E1F2223",
									 -- x"F8F8F8F7", x"F5F4F4F4", x"F7F5F3F2", x"F1F0EEED", x"E6E3DED8", x"D5D5D4D2", x"CBC9C7C7", x"C7C5C4C5",
									 -- x"C2C1BFBE", x"BDBDBEBE", x"C0C0C0C0", x"C1C2C2C2", x"C1C2C2C2", x"C1C1C1C1", x"C1C3C5C5", x"C5C3C3C3",
									 -- x"C1BDB7B3", x"B0ADA9A6", x"A5A19B99", x"99989591", x"928F8E8D", x"8C8A8A8C", x"8C8C8D8D", x"8D8C8B8A",
									 -- x"88888786", x"86868787", x"83868989", x"898B8C8B", x"8B8B8B8A", x"8888898A", x"8A888787", x"8686888B",
									 -- x"8F8C8C8F", x"908E9093", x"93969794", x"94979897", x"9A989695", x"95959595", x"90908F91", x"93949594",
									 -- x"91949696", x"97989897", x"95959596", x"989A9D9E", x"A1A2A5A9", x"AAA9AAAC", x"ACACACB0", x"B6BCC1C3",
									 -- x"C5C3C3C4", x"C3C1C1C2", x"C1C3C4C2", x"C2C3C3C2", x"BFC0B9B4", x"B8BBB8B6", x"AFAFB0B0", x"AFADA8A5",
									 -- x"A5A6A7A6", x"A6A7A5A3", x"9FA0A2A2", x"A2A1A1A0", x"A1A3A4A2", x"A1A09E9C", x"9A979595", x"94919091",
									 -- x"8F8F8E8E", x"8D8E8F90", x"8D8C8B8C", x"8C8B8987", x"88858484", x"84818182", x"84848482", x"81828180",
									 -- x"81818283", x"82818489", x"85888688", x"89888C8A", x"8A8E9191", x"8E8C8C8E", x"93919292", x"8F919594",
									 -- x"92939595", x"96969797", x"98999B9A", x"9897989A", x"9997999E", x"9E9A9899", x"9C9D9FA0", x"A0A1A3A5",
									 -- x"A8A8AAAE", x"AEACABAC", x"A8A6A4A3", x"A5A5A4A3", x"A7A5A29F", x"9C9A9796", x"9795928F", x"8E8E8E8E",
									 -- x"888B8687", x"8C90958F", x"8C898387", x"85828782", x"7D7C7978", x"7878797A", x"78797A7A", x"797A7C7E",
									 -- x"7B7E8286", x"888B8E91", x"908E9195", x"95949493", x"989A9C9E", x"A0A1A09F", x"A4A5A8AB", x"AAA9ACAF",
									 -- x"B5B5B4B0", x"A9A4A5A9", x"ACADACA7", x"A4A29C96", x"90969491", x"94939194", x"969A9998", x"9B9D9EA0",
									 -- x"A0A2A6A8", x"AAA9A49F", x"A3A6ABAF", x"B0AFAEAD", x"B1BABABF", x"C7C7C4BB", x"B4ACADB1", x"AFB0B0AB",
									 -- x"AFAEABA8", x"A8ADB1B2", x"B1B3B2AF", x"ADACA7A1", x"A09C9893", x"91909191", x"8F92979D", x"A4A8A7A3",
									 -- x"9E999899", x"9693918D", x"90929290", x"8F90908F", x"8D8B8885", x"8381807E", x"7E7D7A76", x"726F6F6F",
									 -- x"6C696562", x"615F5C59", x"57535151", x"514F4D4C", x"4C474443", x"423E3B3A", x"3A373637", x"35323030",
									 -- x"2F2B292C", x"2D292728", x"28272626", x"26242220", x"1F1F1F1E", x"1D1C1C1C", x"1F1F1F1F", x"1F202122",
									 -- x"F8F8F7F6", x"F5F4F5F6", x"F6F5F4F3", x"F2F1EFEE", x"E9E5DFD9", x"D6D6D6D4", x"D2CFCBC9", x"C8C6C6C7",
									 -- x"C3C3C2C0", x"BEBEBEBE", x"C1C1C1C1", x"C2C2C3C3", x"C1C2C3C3", x"C2C1C1C1", x"C0C2C4C5", x"C5C4C3C3",
									 -- x"C0BBB4AE", x"ABA7A4A2", x"A4A09B98", x"97959391", x"908E8C8C", x"8A89888A", x"8B8B8C8C", x"8D8D8D8D",
									 -- x"88888786", x"85858585", x"83858788", x"88898988", x"89888887", x"86858586", x"89878584", x"83838588",
									 -- x"8B888889", x"8887898E", x"8F909192", x"92929393", x"93939392", x"92929293", x"91908F8F", x"90919191",
									 -- x"91939596", x"96989999", x"93959797", x"96989DA1", x"A2A3A6A9", x"ABAAABAD", x"AEADAFB4", x"BBC1C5C7",
									 -- x"C8C6C4C3", x"C2C1C1C2", x"C2C3C4C4", x"C5C6C6C4", x"C1C2BCB7", x"BABCB8B6", x"B0B0B1B2", x"B1AEA9A5",
									 -- x"A4A6A6A6", x"A7A8A7A5", x"9EA0A09F", x"A0A2A19D", x"A1A2A2A0", x"9F9E9B97", x"97929193", x"918C8D92",
									 -- x"90908F8E", x"8C8C8E90", x"8B898787", x"89898683", x"857E7C81", x"827E7E81", x"807F7F80", x"7F7D7C7D",
									 -- x"7C7E8080", x"7E7D7F83", x"85838686", x"86888688", x"83888D8E", x"8C8B8D8F", x"8F8C8E8E", x"8C8E9190",
									 -- x"93949596", x"96969797", x"96989997", x"94939496", x"9594969A", x"9B989798", x"9E9E9EA0", x"A4A7AAAB",
									 -- x"B2B1B2B3", x"B3B0ADAB", x"ADABA9A7", x"A7A8A9A9", x"A8A7A6A5", x"A4A19E9C", x"98979591", x"8E8D8F90",
									 -- x"888B8789", x"8D909490", x"898A8886", x"807F8582", x"7E7C7B7A", x"7A7B7C7C", x"7B7E8081", x"81828588",
									 -- x"8385888C", x"8F929394", x"93939397", x"9D9F9EA0", x"A1A09E9E", x"9FA2A6A9", x"ACABABAD", x"AFB1B3B5",
									 -- x"BBBBBAB7", x"B1ADAEB1", x"B8B7B4B2", x"B0ABA49E", x"9A9E9D9C", x"9D99989C", x"9EA2A2A2", x"A6A6A4A4",
									 -- x"A8AAADAF", x"AEA9A7A6", x"A8ACB1B4", x"B4B4B5B6", x"B9BDBFC5", x"C7C7C9C1", x"BAB7B9BB", x"B7B6B6B3",
									 -- x"B5B2ADA9", x"A9ADB1B2", x"B3B5B4B1", x"B0B0ADA8", x"A49F9893", x"9190908F", x"9093999E", x"A4A6A49F",
									 -- x"9A969697", x"94908E89", x"8C8F918E", x"8B8B8B8C", x"89888784", x"82807F7F", x"7B7A7772", x"6D6B6B6C",
									 -- x"6A67625F", x"5E5C5A58", x"55525050", x"504E4B4B", x"4A454141", x"42403C39", x"3A363437", x"342E2D31",
									 -- x"2E2A282B", x"2C2A2726", x"24242424", x"24232220", x"1F212220", x"1D1B1A1A", x"1E1E1F1F", x"1F1F2122",
									 -- x"F4F5F4F4", x"F3F3F4F5", x"F5F4F4F3", x"F2F0EFEE", x"E9E8E4DF", x"DDDBD8D5", x"D7D4D0CC", x"C9C7C6C6",
									 -- x"C4C4C4C2", x"C0BFBFBF", x"C3C3C3C3", x"C3C2C3C3", x"C3C3C4C3", x"C2C1C1C1", x"C1C1C2C2", x"C2C1C1C0",
									 -- x"BEBAB3AC", x"A8A4A09E", x"A09E9B98", x"96959493", x"8D8C8B8C", x"8B898889", x"8989898A", x"8A8B8B8B",
									 -- x"88888685", x"84838382", x"86868584", x"84868788", x"87868585", x"84838485", x"88868585", x"84838487",
									 -- x"87858586", x"8686878A", x"8D8C8D90", x"908D8C8E", x"8C8E9192", x"91909090", x"8F8F8E8E", x"8E8F8F8F",
									 -- x"8E929597", x"989A9998", x"94979897", x"96989DA2", x"A2A3A6A9", x"ABACACAD", x"B0B0B2B8", x"C0C6C9C9",
									 -- x"C9C7C4C2", x"C1C1C1C3", x"C5C3C2C2", x"C4C7C8C8", x"C2C3BFBC", x"BEBCB7B4", x"B3B2B2B4", x"B3AFABA8",
									 -- x"A5A6A6A5", x"A5A7A7A5", x"A2A29F9B", x"9DA2A29D", x"A0A09F9D", x"9C9B9793", x"91909091", x"8F8D8E92",
									 -- x"8F8F8F8D", x"8A8A8B8D", x"89868383", x"8585817D", x"7F7A797B", x"7C7A7B7E", x"7E7C7B7E", x"7D7A797B",
									 -- x"7A7B7D7E", x"7C7B7C7E", x"827D8583", x"84888287", x"81848788", x"88898B8D", x"8A888A8C", x"8B8E908F",
									 -- x"8F909292", x"92929191", x"93969898", x"95939496", x"97959697", x"98989A9D", x"A0A0A1A4", x"A8ADB0B2",
									 -- x"BBBBBBBB", x"B9B6B2B0", x"B3B2B0AE", x"ACACADAE", x"AAABABAB", x"AAA8A4A2", x"9D9B9894", x"91909090",
									 -- x"8A8D8A8E", x"908E908B", x"888B8C88", x"81808480", x"7E80817F", x"7E7F7F7F", x"80838788", x"898B8F93",
									 -- x"94949598", x"9B9C9B9A", x"9EA09C9B", x"A09F9DA1", x"A19F9D9D", x"9EA1A7AB", x"B0AFAFB1", x"B3B5B7B8",
									 -- x"C0C0C0BD", x"B9B7B9BD", x"C4C0BDBB", x"B7B0AAA7", x"A6A7A8A7", x"A5A09FA3", x"A7ABABAA", x"ADABA9AB",
									 -- x"B3B1B1B3", x"B1AEAFB3", x"B1B2B3B3", x"B3B5B8BB", x"BDBFC3CA", x"C8C8CDC6", x"C0C1C2C0", x"BBB7B7B7",
									 -- x"B4B2AFAB", x"A9AAADAF", x"B3B4B4B2", x"B0B0ADAA", x"A6A09994", x"9292918F", x"93979BA0", x"A3A39F9A",
									 -- x"97949596", x"92908F8B", x"878B8D8C", x"8A8A8A8A", x"87868584", x"8281807F", x"78777571", x"6E6B6A69",
									 -- x"6764615E", x"5D5C5A58", x"54525150", x"4E4B4744", x"46444140", x"403E3C39", x"3A373635", x"312D2E32",
									 -- x"302B292A", x"2B292523", x"25242221", x"21212223", x"20222321", x"1D1B1C1E", x"1E1E1E1D", x"1D1E2123",
									 -- x"F1F2F2F2", x"F2F2F3F3", x"F4F4F3F2", x"F1F0F0EF", x"ECEBE9E5", x"E3E1DDD9", x"D7D5D2CF", x"CCCBC9C7",
									 -- x"C6C6C5C4", x"C2C1C1C2", x"C3C4C5C5", x"C4C3C4C5", x"C5C6C5C4", x"C3C1C1C1", x"C2C1C0BF", x"BFBFBFBF",
									 -- x"BDB9B3AD", x"A8A39F9C", x"9B999896", x"9492908F", x"8B8A8A8B", x"8A878686", x"87878787", x"88888888",
									 -- x"88888887", x"87868584", x"86858383", x"83848485", x"85838284", x"84838385", x"84838485", x"84828182",
									 -- x"85838385", x"86868585", x"8987888B", x"8B878687", x"898C8F90", x"8E8D8E90", x"898A8C8E", x"8F909090",
									 -- x"8D919496", x"97999998", x"97979796", x"95979CA0", x"A3A4A7AA", x"ACAFB0B0", x"B4B4B7BC", x"C2C7CACA",
									 -- x"CAC8C5C2", x"C1C1C2C2", x"C4C2C1C2", x"C5C7C8C8", x"C5C5C1BE", x"C0BEB9B8", x"B7B5B4B5", x"B5B1AEAD",
									 -- x"A8A7A5A3", x"A3A5A6A5", x"A3A3A09C", x"9FA5A49F", x"9A9B9A9A", x"9B9B9996", x"90939491", x"90929291",
									 -- x"8B8B8B89", x"87868686", x"86838080", x"81817E7A", x"78797977", x"76767778", x"7B78787A", x"7A777678",
									 -- x"77777879", x"7A7B7A79", x"7C777E7D", x"7E817B81", x"82818081", x"82848585", x"85848789", x"888A8D8B",
									 -- x"8C8E9192", x"91908F8F", x"8F939798", x"97959596", x"9A99999A", x"9A9B9EA1", x"A3A5A8AC", x"AFB3B8BA",
									 -- x"BEC1C3C2", x"C0BDBCBC", x"B7B6B5B3", x"B1AFAEAE", x"B0B0B0AF", x"ADA9A4A1", x"A19E9B99", x"97959390",
									 -- x"8F908D90", x"908C8D89", x"85878C8A", x"85878681", x"7F838582", x"80818486", x"85888C8E", x"9094999D",
									 -- x"9E9E9D9F", x"A1A1A09E", x"A1A6A29E", x"A09D9B9F", x"98999DA2", x"A4A3A4A6", x"B1B3B5B6", x"B6B8BBBD",
									 -- x"C4C5C5C2", x"C0C2C6C9", x"CDCAC7C3", x"BEB8B5B5", x"B1B1B2B2", x"ADAAA9AA", x"AFB3B4B2", x"B2B0B0B6",
									 -- x"BDB9B7B9", x"B9B8B8BB", x"B7B6B4B3", x"B4B6B8B9", x"BDBFC4CD", x"CBCAD0CB", x"CACDCAC4", x"BDB8B7B8",
									 -- x"B6B5B3AF", x"ABABAEB1", x"B3B4B4B2", x"B0AEABA8", x"AAA49C97", x"96969493", x"95999DA0", x"A2A19D98",
									 -- x"96939493", x"9090908C", x"878A8B8A", x"89888785", x"87848180", x"807E7A77", x"77747170", x"6E6B6764",
									 -- x"615F5D5B", x"5A595755", x"51504E4B", x"49464442", x"4242413F", x"3C3A3938", x"37383530", x"2D2F3131",
									 -- x"2E2B2828", x"29272321", x"25242321", x"21212223", x"2021201E", x"1A1A1D20", x"1C1D1E1E", x"1D1E2021",
									 -- x"F1F1F2F2", x"F1F1F1F1", x"F4F4F3F2", x"F1F0F1F1", x"F0EFEBE7", x"E5E4E2DF", x"DBDAD7D3", x"D0CECBC8",
									 -- x"CAC9C7C6", x"C6C5C5C4", x"C3C4C5C6", x"C5C5C6C8", x"C7C8C8C7", x"C5C4C3C3", x"C3C2C0BF", x"BFC0C1C1",
									 -- x"BCB9B4AE", x"A8A39E9B", x"99979593", x"928F8D8B", x"8A89898A", x"88848281", x"85858686", x"86868686",
									 -- x"84858788", x"88878685", x"83828284", x"84828181", x"83807F81", x"82818183", x"82828384", x"83807E7F",
									 -- x"83818082", x"85858280", x"86848588", x"89868586", x"898A8B8A", x"89898C8F", x"87898C8E", x"8F8F8F8F",
									 -- x"90929392", x"93979999", x"9A999897", x"97989C9E", x"A4A6A9AB", x"AFB3B5B4", x"B8B9BBBE", x"C2C5C7C8",
									 -- x"C8C7C4C0", x"BEBEBEBE", x"BFBFC0C4", x"C6C5C5C5", x"C6C5BFBC", x"BDBDBBBC", x"BAB6B4B5", x"B5B1AFAF",
									 -- x"AAA9A6A2", x"A2A3A4A3", x"9FA0A09F", x"A2A5A39E", x"9A9B9A99", x"9A9B9A98", x"90959590", x"8F92918C",
									 -- x"8B8A8988", x"86858382", x"827F7D7D", x"7E7E7C79", x"75787874", x"71727372", x"76747474", x"74737374",
									 -- x"72727172", x"75787876", x"78757879", x"7979777B", x"7E7C7A7C", x"80848584", x"81818586", x"84858887",
									 -- x"8C8F9193", x"94939292", x"8F92979A", x"9A999898", x"9A9B9D9E", x"9E9FA1A3", x"A6ABB0B4", x"B6BABEC2",
									 -- x"C4C8CAC7", x"C4C2C1C1", x"BBBAB8B7", x"B5B2B0AE", x"B2B2B2B1", x"B0ACA8A5", x"A29F9C9A", x"9A989592",
									 -- x"92918B8E", x"8D898C8B", x"88858A89", x"87898480", x"83878884", x"82868B8D", x"8B8D9195", x"989DA1A4",
									 -- x"A09F9FA0", x"A2A3A2A1", x"A0A3A3A0", x"9F9E9D9F", x"99999CA1", x"A3A3A5A9", x"AEB3B6B6", x"B6B8BCBF",
									 -- x"C5C6C6C4", x"C4C7CCCF", x"CDCDCBC7", x"C3BFBDBD", x"B8B8BAB9", x"B4B3B3AE", x"B3B8BAB8", x"B7B4B5BC",
									 -- x"C1BFBFC1", x"C3C2BEBC", x"B7B6B4B4", x"B5B5B5B4", x"B3B7BBC6", x"C7C4CAC8", x"CED1CCC3", x"BFB9B6B9",
									 -- x"B8B6B3B0", x"ADACAFB4", x"B3B4B3B1", x"AEABA8A7", x"AAA59E99", x"97969594", x"979A9D9F", x"A0A09D99",
									 -- x"96949491", x"8D8D8E8A", x"898B8A88", x"8684827F", x"83817E7E", x"7E7D7874", x"7673706F", x"6E6B6560",
									 -- x"5E5C5B59", x"58565553", x"504F4B47", x"45464746", x"4042423F", x"3B393838", x"3336332C", x"2B303230",
									 -- x"2C2A2929", x"29272524", x"23242424", x"23222121", x"22211F1C", x"191A1D20", x"191C2020", x"1F1E1D1E",
									 -- x"F0F0F0EF", x"EFEFF0F1", x"F3F3F2F1", x"EFEFF0F2", x"F1F0ECE8", x"E6E6E5E2", x"E0DFDCD7", x"D4D3D0CC",
									 -- x"D0CDCAC8", x"C9C9C8C6", x"C3C5C6C7", x"C6C6C7C9", x"C7C9CBCB", x"CAC8C6C5", x"C4C2C0BF", x"C0C1C1C1",
									 -- x"BCB9B4AD", x"A7A19D9A", x"99979391", x"908E8C8A", x"8B898888", x"86838181", x"82838484", x"85848483",
									 -- x"81828586", x"86858382", x"817F7F82", x"82807E7E", x"807C7B7E", x"7F7C7C7F", x"7F7F8182", x"817F7E7E",
									 -- x"7F7F7F80", x"81828180", x"84848486", x"87878685", x"85868686", x"85858788", x"87898B8D", x"8D8D8D8E",
									 -- x"91929291", x"92959798", x"9A999997", x"97989B9E", x"A4A6A9AC", x"B1B7B9B8", x"BCBDBFC0", x"C1C2C4C5",
									 -- x"C2C3C0BD", x"BBBBBBB9", x"BBBBBDC1", x"C2C0C1C2", x"C5C4BFBC", x"BDBBB9BA", x"BAB5B3B5", x"B4B0AEAF",
									 -- x"ABAAA7A4", x"A3A4A3A2", x"A09F9FA0", x"A2A29F9D", x"9C9D9C99", x"97989897", x"9293918E", x"8D8E8D8A",
									 -- x"8D8B8886", x"86858381", x"7F7D7B7A", x"7A7A7977", x"75757474", x"726F6E6E", x"7272716E", x"6E6F7070",
									 -- x"6E6F6E6D", x"6F727473", x"77767378", x"78737677", x"7877787B", x"7F838585", x"80818688", x"84858889",
									 -- x"8A8C8E90", x"92939495", x"96989C9F", x"A0A09E9D", x"9EA0A2A2", x"A3A5A8AA", x"AEB2B8BC", x"BFC3C8CC",
									 -- x"CED0D0CC", x"C9C8C6C5", x"C3C1BEBD", x"BCBAB7B4", x"B3B4B4B4", x"B4B2AFAD", x"A5A3A09E", x"9C9A9896",
									 -- x"94928C8F", x"8E898C8D", x"90888C8B", x"898C8786", x"8D908F8C", x"8D909291", x"9294979B", x"9FA2A3A4",
									 -- x"A5A5A5A5", x"A6A7A8A8", x"A8A8A8A4", x"9E9B9893", x"9D9A9A9C", x"9E9FA6AE", x"A9AEB2B3", x"B4B8BCBF",
									 -- x"C4C7C8C6", x"C6CACDCE", x"CBCECECB", x"C8C6C2BD", x"BDBCBFBD", x"B9BDBDB3", x"B6BBBEBF", x"BFBBBABF",
									 -- x"BFC1C3C6", x"C7C6C1BB", x"B6B6B4B2", x"B1B0B1B1", x"ABB0B1BA", x"BFBBBEC0", x"C7CBC6BF", x"BFBCB9BB",
									 -- x"B7B3B0B0", x"B0AFAFB0", x"B0AFAEAB", x"A7A5A4A5", x"A3A09B97", x"94949494", x"999C9E9F", x"9F9F9C99",
									 -- x"97959591", x"8C8C8D89", x"87898A86", x"82807F7E", x"807F7E7D", x"7D7B7774", x"72706D6B", x"6A66615E",
									 -- x"5E5C5957", x"55535352", x"4F4F4D48", x"46464746", x"3F41413E", x"3C3B3937", x"3535332F", x"2E2F2F2C",
									 -- x"2A2A2B2A", x"29282727", x"22232424", x"23222122", x"2221201E", x"1C1D1E20", x"1A1D1F1F", x"1D1C1D1E",
									 -- x"EEEEEDEC", x"EDEEF0F2", x"F1F1F0EF", x"EDEDEFF1", x"F0EFECE9", x"E8E7E5E1", x"DFDFDDD9", x"D8D9D8D5",
									 -- x"D5D0CCCA", x"CBCCCAC7", x"C5C7C8C7", x"C6C5C7C8", x"C7C9CDCE", x"CECBC8C6", x"C4C2C1C0", x"C0C0BFBE",
									 -- x"BDB9B3AC", x"A5A09C9A", x"9894908E", x"8D8D8B89", x"8B898887", x"86848385", x"7F808183", x"83838281",
									 -- x"81828586", x"8684807E", x"827E7C7E", x"7F7E7E7F", x"7E7A787B", x"7C79797B", x"7B7B7D7F", x"7F7D7D7E",
									 -- x"7C7D7E7E", x"7F818283", x"82838383", x"84858481", x"7F828486", x"85848280", x"8486898A", x"8C8D9091",
									 -- x"8F919393", x"93959695", x"96979796", x"9494989C", x"A3A5A8AB", x"B1B8BAB9", x"BEBFC1C1", x"BFBFC1C3",
									 -- x"BFC0BFBD", x"BBBCBCBA", x"B9B8B9BB", x"BBBBBDC1", x"C6C7C4C2", x"C2BDB7B6", x"B8B4B2B4", x"B4AFADAE",
									 -- x"AAAAA8A6", x"A4A4A3A1", x"A6A3A1A1", x"A19F9E9F", x"9B9C9B98", x"95969798", x"94918E8E", x"8F8E8D8D",
									 -- x"8D8A8583", x"8483817F", x"7E7D7B79", x"78777675", x"77727074", x"746E6B6D", x"6F716F6B", x"6B6E6F6E",
									 -- x"6E706F6C", x"6B6E7070", x"74756F76", x"76707675", x"7677787A", x"7C7D7E7E", x"8083898B", x"87888C8E",
									 -- x"8E8F9194", x"96999C9D", x"9FA0A1A4", x"A7A7A5A3", x"A7A8A8A7", x"A8ACB2B6", x"B8BBBFC4", x"C8CDD3D6",
									 -- x"D5D5D4D2", x"D1D2D0CD", x"CBC8C5C3", x"C3C2BEBB", x"BAB9B9B8", x"B7B5B2B0", x"ABAAA7A3", x"9F9D9C9C",
									 -- x"98969296", x"958E9090", x"978B908F", x"90949195", x"95989897", x"999B9790", x"999A9DA0", x"A4A4A2A0",
									 -- x"A4A4A4A4", x"A4A5A6A7", x"A6A3A6A5", x"A0A09D94", x"9998999D", x"9E9EA3AA", x"A8ACAFB0", x"B3B9BEC0",
									 -- x"C6C9CBCA", x"CACCCECE", x"CDD2D3D0", x"D0CFC7BD", x"C1C1C4C2", x"BFC5C6B9", x"BABFC2C6", x"C8C3BFC2",
									 -- x"BCC0C4C5", x"C6C6C2BB", x"B7B6B3AF", x"ABAAACAF", x"ACB1AEB6", x"BDB7B8BD", x"BFC4BFBB", x"C0C0BDBF",
									 -- x"B4B0AEB2", x"B5B3AEAB", x"ACAAA7A4", x"A19FA1A3", x"9E9C9995", x"94949596", x"9C9E9F9F", x"9E9D9B98",
									 -- x"97969692", x"8D8D8E8A", x"81868884", x"7F7D7E80", x"8180807D", x"7A75726F", x"6A696866", x"63605E5C",
									 -- x"5D5B5754", x"51505050", x"4D4F4E4A", x"4644423E", x"3D3E3D3B", x"3A3A3834", x"3A363433", x"322E2B29",
									 -- x"28292A29", x"27262525", x"24242322", x"20212324", x"1F1F1E1E", x"1E1E1E1E", x"1E1F1E1C", x"191A1E21",
									 -- x"ECECECEC", x"ECEDEEF0", x"F1EFECEC", x"EEEFEFEF", x"EFEEEDEB", x"EAE8E5E4", x"DFDEDDDE", x"E0E0DEDC",
									 -- x"DAD9D8D5", x"D1CFCDCD", x"CCCAC9C8", x"C9C9C8C7", x"C8CACBCD", x"CDCDCCCB", x"C5C2BFBF", x"BFBEBDBD",
									 -- x"BDB7AFAA", x"A6A29D98", x"9A969391", x"8F8C8989", x"88878686", x"8887837F", x"7F808080", x"7F808284",
									 -- x"84838381", x"80808182", x"7E7E7E7D", x"7D7E7D7A", x"7A797979", x"7876787A", x"7A7C7C7B", x"79797B7D",
									 -- x"7D7E7E7B", x"7B81827A", x"807F7E7F", x"80807E7C", x"837F7D81", x"82807E80", x"83858789", x"8B8D8F90",
									 -- x"8B8F9394", x"95979796", x"96999997", x"95969695", x"9EA0A1A6", x"AFB3B7BE", x"BCC0BFBD", x"C1C2C0C0",
									 -- x"BEBEBDBB", x"BAB9B8B6", x"B8B8B9B9", x"BBBDBDBC", x"C4C2C1C1", x"BDB7B6B8", x"B1B0AEAD", x"AEB1AFAB",
									 -- x"A8A7A5A4", x"A3A4A3A3", x"A0A1A19F", x"9EA09F9D", x"9A989797", x"97969390", x"95918E8F", x"908E8C8A",
									 -- x"88858384", x"83807E7F", x"847C7576", x"7977736F", x"72726F6D", x"6E706E6B", x"6E6D6A67", x"67696969",
									 -- x"6A69696A", x"6A6A6C6F", x"6F6F7072", x"74747372", x"76787776", x"76797C7C", x"83888A8B", x"8D8D8E93",
									 -- x"96969698", x"9A9EA1A3", x"A7A5A7AB", x"ADACACAD", x"A8ACB0B1", x"B2B6B9BB", x"BEC1C7CB", x"CFD4D8DC",
									 -- x"DBDCD8D1", x"CED2D5D5", x"D6D1CAC7", x"C6C6C5C2", x"C1BFBDBC", x"B8B5B5B7", x"B3AEA9A7", x"A39E9B9B",
									 -- x"98969495", x"9796938F", x"94939091", x"9696969A", x"9CA09E9C", x"9FA09E9E", x"9EA1A5A9", x"ABA6A3A7",
									 -- x"AAA6A4A6", x"A6A3A4A8", x"A6A4A3A5", x"A5A29A94", x"969A9799", x"9A9CA3A1", x"A8A6A9B0", x"B3B2B6BC",
									 -- x"BABCC1C6", x"C7C7CACE", x"C8C9CDD4", x"D3CBC3C0", x"C2C4C3C1", x"C4C9C9C6", x"C1C1C4C9", x"CAC9C6C6",
									 -- x"C2C2C6CA", x"C8C0B9B7", x"B7B3B1B1", x"B0ADACAE", x"B1B5B7B6", x"B5B6B7B7", x"BEBCC0C5", x"C0BCBCBC",
									 -- x"B7AFAAAD", x"B2B0A8A2", x"AAA6A4A4", x"A4A09A96", x"97969793", x"8C8E9699", x"9D9C9998", x"98989898",
									 -- x"95989792", x"8D8C8C8C", x"82848382", x"85848181", x"80807E78", x"726F6F71", x"6A696765", x"64615C58",
									 -- x"53555554", x"5352504D", x"4A494949", x"4845413E", x"3C3C3B3A", x"39373635", x"33333231", x"302E2C2A",
									 -- x"2B282424", x"272A2722", x"23242423", x"22222222", x"201D1B1D", x"1E1D1D1D", x"1D1C1B1B", x"1C1E2022",
									 -- x"ECECECEC", x"EBEAEBEB", x"EEEEEDED", x"ECEDEEEE", x"EDEDECEB", x"EAE9E7E5", x"E2E1E1E2", x"E3E4E2E0",
									 -- x"DFDEDEDC", x"D9D6D3D1", x"D3D2CFCD", x"CCCBCAC9", x"CACBCBCC", x"CCCDCDCC", x"C9C5C2C1", x"BFBCBAB9",
									 -- x"B4B0ABA7", x"A39F9B98", x"9693908F", x"8E8C8A8A", x"86858586", x"87878482", x"7E7F7F7E", x"7E7E7F80",
									 -- x"7D7F8182", x"817F7E7D", x"81817F7C", x"7B7B7977", x"79787878", x"77767779", x"78797A7A", x"79797B7C",
									 -- x"7C7A7B7A", x"7A7F807B", x"82817F7F", x"7F7E7C7A", x"7A7A7C7E", x"7C797C81", x"82848789", x"8A8C8E90",
									 -- x"8F90908F", x"91949493", x"95979896", x"94959695", x"9C9FA0A3", x"A9ADB2BA", x"BCC0BFBE", x"C1C1BEBE",
									 -- x"BCBCBBBA", x"B9B8B7B6", x"B4B5B5B6", x"B7B9BBBB", x"C2C1C0BF", x"BDB8B5B4", x"B2B1AEAC", x"ACADACA9",
									 -- x"A6A6A5A4", x"A4A4A3A2", x"A1A2A2A0", x"9F9F9D9B", x"97969697", x"98979492", x"95908D8D", x"8D8C8A89",
									 -- x"85838383", x"827F7E80", x"77767676", x"74717173", x"6E6D6C6B", x"6E706D68", x"6A696968", x"68686868",
									 -- x"6465686B", x"6B69696A", x"70707072", x"74767777", x"76797A7B", x"7D808384", x"858B8D8F", x"92929296",
									 -- x"98999B9D", x"A0A3A6A8", x"ACADB0B3", x"B4B3B4B6", x"B4B7B9B9", x"B9BDC0C1", x"C3C6CACE", x"D2D7DDE0",
									 -- x"DDDFDCD5", x"D2D5D8D8", x"DAD5D0CD", x"CCCCC9C7", x"C2C0BEBD", x"BBB8B8B9", x"B7B2ADAB", x"A8A3A09F",
									 -- x"9B9A9897", x"96959493", x"96969496", x"9B9D9DA1", x"A0A6A6A4", x"A5A4A3A4", x"A6A9AAAA", x"AAA6A4A8",
									 -- x"A6A8A9A9", x"AAAAA9A8", x"A7A6A5A4", x"A2A09C99", x"989A989D", x"9E9DA19F", x"A6A5A8AD", x"B1B1B2B6",
									 -- x"B3B4B7BB", x"BDC0C8CF", x"CBC7C8CC", x"CEC9C3C2", x"BEBFBFC2", x"C8CFD2D1", x"CACACBCD", x"CCC8C3C1",
									 -- x"BEC1C3C2", x"BFBBB7B4", x"ADAEB0B1", x"AFACABAC", x"ACAFB1B1", x"B1B3B5B6", x"BCBBBEBE", x"BBBBBDBA",
									 -- x"B5B0ACAD", x"AEACA7A4", x"ABA7A3A2", x"A19C9693", x"93949797", x"92939798", x"9A989695", x"94949393",
									 -- x"91918E8A", x"88888684", x"8283807F", x"82807C7B", x"7C7A7773", x"6F6C6B6B", x"6866625F", x"5D5D5C5A",
									 -- x"54555552", x"514F4D4A", x"4A484645", x"4442403E", x"3D3D3C3B", x"39373534", x"33312F2E", x"2D2E2E2E",
									 -- x"2A2A2827", x"28282623", x"25262625", x"23222121", x"1F1E1E1F", x"1F1E1F21", x"201E1D1D", x"1F212323",
									 -- x"EAEBEBEA", x"E9E8E8E8", x"EAECEEED", x"ECEBECED", x"ECEBEBEB", x"EAE9E8E6", x"E4E3E3E4", x"E5E6E5E3",
									 -- x"E4E4E3E3", x"E2DFDAD7", x"D9D7D5D1", x"CECCCBCB", x"CCCCCCCB", x"CCCDCDCE", x"CAC6C3C1", x"BEBAB6B4",
									 -- x"AFAEABA7", x"A39F9C9A", x"96928F8E", x"8C8A8787", x"84848383", x"84838281", x"7D7D7C7C", x"7D7C7C7B",
									 -- x"787B7E7F", x"7F7D7B7A", x"7C7C7B79", x"797A7978", x"78777778", x"76757577", x"77777878", x"79797979",
									 -- x"7B777779", x"787A7C7A", x"7E7E7E7F", x"7F7C7976", x"78787A7C", x"7A787C81", x"82848789", x"898A8D8F",
									 -- x"91908E8D", x"8F929291", x"93959695", x"94959696", x"9DA0A1A3", x"A6A8AEB7", x"B6BABABA", x"BDBCBABA",
									 -- x"B9B8B8B7", x"B7B6B6B6", x"B3B4B4B4", x"B4B4B6B8", x"BABABABB", x"BBBBB7B3", x"B1B0AEAB", x"A9A9A9A8",
									 -- x"A3A2A2A2", x"A2A1A09F", x"9FA0A1A0", x"9E9D9B98", x"95949495", x"96959391", x"928E8B8A", x"8B898888",
									 -- x"84838282", x"7F7D7C7C", x"76777978", x"74707073", x"6E6E6D6D", x"6F706C67", x"6666676A", x"69666668",
									 -- x"6A686767", x"67676A6D", x"6E6E6E70", x"7376797B", x"787B7E7F", x"82868888", x"898E9194", x"98989799",
									 -- x"9C9EA1A4", x"A6A9ACAE", x"B2B5BABD", x"BCBBBCC0", x"C0C2C3C1", x"C1C4C6C8", x"CACBCED1", x"D5DAE0E3",
									 -- x"E1E3E0DB", x"D8DADDDD", x"DDD9D4D1", x"D1D0CECB", x"C6C2C0BF", x"BFBEBDBE", x"BBB6B1AF", x"ADAAA7A4",
									 -- x"9F9F9D9A", x"96959698", x"9B9C9A9C", x"A1A3A3A8", x"A4ABACAA", x"A9A7A6A9", x"A9ADACA9", x"AAA9A9AB",
									 -- x"A5AAABA9", x"A9ACAAA5", x"A6A6A4A1", x"9F9E9D9E", x"9A9A979D", x"9F9B9F9F", x"A6A6A8AB", x"AFB1B1B1",
									 -- x"B1B2B5B7", x"BABFC9D1", x"D0CBC8CC", x"CECBC7C5", x"C0BDBEC5", x"CDD3D7D8", x"D7D5D5D4", x"D1CBC5C2",
									 -- x"BCC0C0BA", x"B7B7B5B1", x"AAAEB1B0", x"AEADADAD", x"ACAEAFAE", x"AEB1B4B6", x"B5B6B8B6", x"B4B8B8B1",
									 -- x"B3B0ADAB", x"A9A6A3A3", x"A5A09D9D", x"9D9A9795", x"93929596", x"93939695", x"94939292", x"9191908F",
									 -- x"8F8D8886", x"8686837F", x"80817E7D", x"7F7C7776", x"7674716F", x"6D6B6967", x"65625E5B", x"58575858",
									 -- x"5353514E", x"4C4C4A47", x"47454342", x"41403E3D", x"3D3D3D3C", x"3A383534", x"3634302E", x"2D2D2D2D",
									 -- x"282A2B29", x"27262524", x"25252625", x"23222121", x"1F1F2020", x"1F1E1F22", x"211F1D1D", x"1F212223",
									 -- x"E9E9E9E8", x"E7E7E7E8", x"E8EAECED", x"ECEBEBEB", x"EBEAEAEA", x"EAE9E8E7", x"E5E5E5E5", x"E6E7E6E6",
									 -- x"E7E6E5E6", x"E6E3DEDB", x"D9D8D6D2", x"CECCCCCD", x"CDCDCCCC", x"CCCCCDCE", x"C8C5C2C0", x"BEB9B5B3",
									 -- x"B1AFACA9", x"A6A29E9B", x"96928F8D", x"8B888585", x"82828180", x"7F7E7D7D", x"7C7B7A7A", x"7B7B7977",
									 -- x"7778797A", x"79797A7A", x"76767574", x"75777877", x"78777677", x"76747475", x"77777777", x"78787776",
									 -- x"7A757579", x"77767776", x"77787A7D", x"7D7B7773", x"7B78777A", x"7C7C7D7E", x"81848889", x"89898C8E",
									 -- x"8D8D8D8D", x"8E8F8F8E", x"91939494", x"94949697", x"9EA1A2A3", x"A7A7ABB2", x"AFB3B3B4", x"B7B7B6B8",
									 -- x"B7B6B5B5", x"B5B4B5B6", x"B3B3B4B3", x"B0AEAFB1", x"B2B5B6B5", x"B6B9B7B2", x"AEAEADAB", x"A8A7A7A7",
									 -- x"A1A09F9F", x"9F9E9C9C", x"9A9B9C9B", x"9B9A9998", x"95949392", x"91908E8D", x"8F8C8989", x"8A888787",
									 -- x"8683817F", x"7D7B7876", x"7B787676", x"76757370", x"70706F6F", x"6E6C6966", x"6565676B", x"69656569",
									 -- x"6F6B6867", x"66676B6F", x"6C6E7072", x"75787C7E", x"7F828484", x"86898B8B", x"9094979A", x"9F9F9D9F",
									 -- x"A3A5A9AB", x"AEB2B6B8", x"BCC0C4C6", x"C5C4C5C7", x"CACBCCCA", x"CACCCDCD", x"CFD0D2D5", x"D9DDE1E3",
									 -- x"E6E6E5E0", x"DEDFE0E1", x"DDD9D5D2", x"D2D2D1CF", x"CBC7C3C2", x"C3C4C2C1", x"BCB8B4B2", x"B2B0ADAA",
									 -- x"A5A4A19E", x"9B999A9C", x"A1A1A0A1", x"A5A5A5AA", x"A8ADADAB", x"AAA8A7AB", x"ACB1AEAA", x"ABADACAD",
									 -- x"ACAEAEAA", x"A8AAA9A5", x"A5A4A2A0", x"9E9D9D9D", x"9A99959A", x"9A959CA0", x"A3A5A6A7", x"ACB1B2AE",
									 -- x"B0B3B7BA", x"BCC1C8CE", x"CECBCACC", x"CDCAC6C4", x"C1BCBDC7", x"D0D5D9DD", x"DDDAD8D7", x"D4CECAC8",
									 -- x"BFBEBBB7", x"B4B2B1AF", x"AEB0AFAC", x"ABADAFAF", x"AFAFAEAD", x"ACAFB2B4", x"AEAFB2B3", x"B1B2B0A9",
									 -- x"B0AEABA8", x"A5A2A09F", x"9E9A9798", x"99989796", x"96929191", x"8F8F9291", x"8D8D8C8C", x"8D8C8B8A",
									 -- x"8D898584", x"8585827F", x"7C7E7C7A", x"7B777474", x"706F6E6C", x"6B696664", x"61605E5C", x"58545253",
									 -- x"52514E4C", x"4B4B4A48", x"42424243", x"43413E3B", x"3D3D3D3C", x"3B383534", x"38363331", x"2F2D2B29",
									 -- x"282A2B29", x"26262524", x"22232424", x"23222121", x"21202021", x"1F1D1E20", x"1D1D1D1D", x"1C1D2021",
									 -- x"EBEAE9E7", x"E5E6E7E8", x"E8E8E9EB", x"EDEDECEA", x"EAEAEAEA", x"E9E9E7E6", x"E7E7E6E7", x"E7E8E8E7",
									 -- x"E7E6E5E5", x"E6E4E1DD", x"DBDAD8D4", x"D0CFCFD0", x"CECECDCD", x"CDCCCCCC", x"C7C4C2C1", x"BFBBB7B5",
									 -- x"B4B0ACA9", x"A7A49E9A", x"93908D8C", x"8B898787", x"80807F7D", x"7C7B7B7A", x"7A797979", x"7A797674",
									 -- x"76777777", x"7677787A", x"76767472", x"72737371", x"74727274", x"74737374", x"76767676", x"76757371",
									 -- x"76717377", x"75737473", x"75767779", x"7A797877", x"79777679", x"7B7D7D7D", x"81838788", x"89898B8D",
									 -- x"898A8B8B", x"89898B8E", x"8F909293", x"93949698", x"9B9E9EA1", x"A6A6A6AA", x"ACAFAFB0", x"B3B3B3B7",
									 -- x"B5B4B3B5", x"B5B3B3B5", x"B2B2B2B2", x"AEAAAAAC", x"B1B4B4B1", x"AFB0B0AE", x"ABACADAC", x"A9A5A4A5",
									 -- x"A29F9D9D", x"9D9A9A9B", x"98989797", x"97969797", x"9694928F", x"8E8D8C8B", x"8D8B8989", x"88868484",
									 -- x"83807C7B", x"7C7B7774", x"76726F70", x"73767471", x"6F6F6F6D", x"69666566", x"6767696B", x"69666669",
									 -- x"6969696B", x"6B6A6B6D", x"6F72777A", x"7C7E8183", x"87898B8B", x"8C909393", x"999EA0A2", x"A6A6A6A9",
									 -- x"AEB0B2B5", x"B8BCC1C5", x"CACCCFD0", x"CFCFCFCF", x"D2D4D5D4", x"D4D4D4D3", x"D2D3D5DA", x"DFE3E4E5",
									 -- x"E9E9E7E4", x"E1E1E2E3", x"DEDBD7D5", x"D5D5D5D4", x"D2CDC8C5", x"C6C6C3C0", x"C0BDB9B7", x"B6B5B2AF",
									 -- x"AAA7A4A2", x"A1A09F9E", x"A2A4A2A4", x"A8A8A8AD", x"AEAFACAA", x"ACABAAAD", x"AEB3B0AC", x"ADAFADAD",
									 -- x"B5B4B3B2", x"AFADAAA9", x"A6A5A2A1", x"9F9D9A98", x"97979499", x"97929AA0", x"9FA1A2A2", x"A7AEB0AD",
									 -- x"ADB1B5B8", x"BBBFC4C7", x"C5C5C5C6", x"C6C4C2C2", x"BDB9BCC8", x"D3D8DCE1", x"DDDAD7D6", x"D4D1CFCE",
									 -- x"C5BEB8B8", x"B6B0ACAD", x"B0AFABA8", x"A9ABACAC", x"AEACAAA9", x"A9AAADAF", x"B0ACAEB2", x"B0ADACA8",
									 -- x"ABAAA7A5", x"A4A29F9C", x"9D999595", x"95949494", x"98918F8F", x"8D8C8E8D", x"88878787", x"86858482",
									 -- x"8482807F", x"7F7E7D7C", x"777B7A77", x"75716F72", x"6A6B6B69", x"66636160", x"5F5E5D5D", x"59545151",
									 -- x"52514E4B", x"4B4D4C49", x"42424243", x"4342403D", x"3C3C3D3C", x"3B383634", x"36343231", x"2F2E2C2B",
									 -- x"2A2A2927", x"27282725", x"23242424", x"23222222", x"23201F20", x"211F1E1E", x"1C1F201E", x"1C1B1F22",
									 -- x"EDECEAE7", x"E6E5E6E7", x"E8E7E8EA", x"ECEDEBE9", x"EAE9E9E9", x"E8E7E6E5", x"E5E5E5E5", x"E5E5E5E5",
									 -- x"E7E6E5E5", x"E5E4E2E0", x"DFDEDBD8", x"D5D3D3D3", x"CFCFCFCF", x"CECDCBCA", x"C9C6C4C4", x"C2BFBBBA",
									 -- x"B8B3ADA9", x"A8A59F9B", x"94918D8C", x"8A878584", x"7F7E7D7C", x"7B7B7A79", x"77777778", x"78777574",
									 -- x"73757677", x"77777676", x"77767572", x"7172716F", x"6D6C6C6F", x"70706F70", x"73737373", x"72706F6E",
									 -- x"6F6C6F73", x"71707171", x"77767574", x"7576787A", x"7376797A", x"7A7A7D81", x"7E808385", x"8788898A",
									 -- x"8C8C8C8A", x"87868B91", x"8E8E9092", x"93939597", x"989A9B9F", x"A5A4A3A6", x"AAACABAB", x"ADACADB2",
									 -- x"B3B1B2B4", x"B5B2B2B4", x"B5B3B3B3", x"B0ACABAE", x"ADAFAFAC", x"AAAAACAD", x"ABABACAC", x"A8A4A1A1",
									 -- x"A39F9D9D", x"9C99999A", x"99979695", x"94939394", x"9392908E", x"8C8C8C8C", x"8C8A8887", x"85828080",
									 -- x"7D7B7978", x"7A7B7874", x"7172716F", x"6E707171", x"6F6E6E6C", x"6967676A", x"696B6C6C", x"6B69696A",
									 -- x"6A6A6B6E", x"6F707376", x"757A7F81", x"82838688", x"8B8D9091", x"94999C9D", x"A1A6A9AA", x"ADADADB1",
									 -- x"B7B9BCBE", x"C0C5CACF", x"D6D8D9D8", x"D8D8D8D7", x"D9DBDCDB", x"DADAD9D6", x"D5D6DAE0", x"E6EAEBEA",
									 -- x"ECEBE9E6", x"E3E2E3E4", x"E2E0DDDB", x"DBDCDBDB", x"D7D3CDC8", x"C7C6C3C0", x"C6C4C1BE", x"BCBAB7B4",
									 -- x"B1ADA9A8", x"A8A8A5A2", x"A4A6A6A8", x"ACACADB3", x"B1B1ADAB", x"AEADACB0", x"ACB0AEAD", x"B0B1B0B1",
									 -- x"B9B9B9B9", x"B6B1ACAB", x"AAA8A5A3", x"A19D9995", x"9597969A", x"9893999C", x"9C9EA0A1", x"A6ACADAC",
									 -- x"ADB0B4B7", x"BBC1C5C6", x"C2C2C1C0", x"C0C0C3C5", x"BDBBC0CB", x"D4D8DCE0", x"DDDAD8D7", x"D5D3D2D3",
									 -- x"CCC2BDBE", x"BBB2ADAF", x"AFABA9AA", x"ABABAAA9", x"ABA9A8A8", x"A8A9ABAD", x"B1AAAAAD", x"AAA8A9AA",
									 -- x"A6A5A4A3", x"A3A4A19E", x"9D999594", x"94939394", x"958F8E90", x"8D8B8A88", x"86858483", x"82817F7D",
									 -- x"7D7B7A79", x"78767677", x"73777571", x"6E6A686C", x"69696967", x"635F5D5C", x"5E5B5959", x"57545354",
									 -- x"514F4C49", x"494B4A47", x"46444241", x"42424140", x"3D3D3D3C", x"3B393736", x"3835312E", x"2D2C2C2B",
									 -- x"2E2C2A28", x"2A2B2A26", x"27272625", x"24232323", x"23212021", x"23222020", x"1F222422", x"1F1E2125",
									 -- x"ECECEBE9", x"E7E6E6E7", x"E7E7E8E8", x"E9E9E9E9", x"E8E8E8E8", x"E8E7E5E4", x"E3E3E3E2", x"E1E1E2E3",
									 -- x"E4E4E5E4", x"E4E3E1E1", x"E0DEDCDA", x"D8D7D5D5", x"D2D2D2D1", x"CFCDCCCB", x"C9C6C5C5", x"C5C2C0BF",
									 -- x"BEB9B1AB", x"A7A39F9C", x"97928E8C", x"89858281", x"807D7B7B", x"7B7A7876", x"74757676", x"75757475",
									 -- x"72747677", x"77767574", x"75757471", x"7171706E", x"6C6A6A6C", x"6D6C6B6B", x"6C6E6F6E", x"6C6B6B6C",
									 -- x"6A686A6C", x"6A6C6E6E", x"71707070", x"71727475", x"70747879", x"78787B7D", x"7B7C7E81", x"84868685",
									 -- x"8C8B8A89", x"87878B90", x"8C8C8E91", x"91919396", x"94989A9E", x"A3A3A3A8", x"A5A8A7A8", x"AAA8A8AE",
									 -- x"B0AEB0B4", x"B5B2B2B4", x"B8B4B2B2", x"B1AEAEB1", x"ABA9A8A8", x"A8A8A9AB", x"AAA9A9AA", x"A7A29F9F",
									 -- x"A19D9B9C", x"9B989799", x"97959494", x"92908F90", x"8D8D8D8C", x"8B8B8B8B", x"8A868382", x"807E7D7E",
									 -- x"7B7C7A77", x"76767573", x"72757572", x"6F6F7071", x"72706E6F", x"6E6D6C6E", x"6B6E6F6D", x"6D6F6E6A",
									 -- x"71707073", x"76797E83", x"7F838686", x"85878B8F", x"90939699", x"9CA1A4A5", x"A7AFB3B5", x"B7B6B6BB",
									 -- x"C0C3C6C9", x"CBCFD4D8", x"DFE3E4E2", x"DFDFE1E1", x"E2E3E2E0", x"DFDEDCD9", x"DBDCDFE5", x"EBEFEFED",
									 -- x"EEECEAE6", x"E3E2E3E5", x"E6E5E3E2", x"E2E1DFDE", x"DAD7D2CC", x"CACAC8C4", x"C8C9C7C3", x"C0BFBDBA",
									 -- x"BCB7B3B1", x"B1B0ADAA", x"ABADADAF", x"B2B1B2B7", x"B4B4B2B1", x"B2B0B0B5", x"B3B4B3B3", x"B7B6B4B8",
									 -- x"BCBEBDB9", x"B6B3AFAA", x"AAA9A6A3", x"9F9C9998", x"97999597", x"97959997", x"9A9C9FA2", x"A5A8A9A9",
									 -- x"ACAFB3B7", x"BEC4C6C4", x"C3C2BFBD", x"BEC0C3C5", x"C2C4C9D1", x"D6D8DADC", x"DBD9D7D7", x"D6D4D3D3",
									 -- x"CCC7C3C1", x"BCB3B0B2", x"ADA8A7AB", x"ACA7A6A8", x"ABA9A8A9", x"AAA9ABAD", x"ADA9A9A9", x"A5A5A8A8",
									 -- x"A4A4A3A2", x"A2A4A4A1", x"A09C9896", x"95939394", x"908A8B8D", x"89858382", x"8281807F", x"7E7D7C7A",
									 -- x"7A777676", x"74717172", x"71726E6B", x"6A676668", x"66656464", x"62605D5B", x"5B565455", x"55535355",
									 -- x"4D4C4947", x"484B4A47", x"47454241", x"4141403F", x"3F3F3E3D", x"3B3A3837", x"39363330", x"2E2D2C2C",
									 -- x"2E2E2C2A", x"2B2C2A26", x"28282725", x"24232424", x"22212122", x"22212020", x"23242423", x"22212325",
									 -- x"E9EAEAEA", x"E9E8E7E7", x"E7E8E8E8", x"E6E6E7E8", x"E7E7E7E7", x"E7E7E5E4", x"E4E4E4E3", x"E2E1E2E3",
									 -- x"E2E3E4E4", x"E3E2E1E0", x"DDDCD9D8", x"D8D8D6D4", x"D5D4D3D1", x"D0CECCCB", x"C7C4C4C5", x"C6C4C3C2",
									 -- x"C1BCB4AC", x"A59F9C9A", x"94908C8B", x"89858382", x"807D7A79", x"79787571", x"72737575", x"74737475",
									 -- x"73747575", x"75757575", x"75757471", x"6F6F6D6A", x"6E6C6B6C", x"6B696766", x"67696B6A", x"6968696B",
									 -- x"68666767", x"64676B6A", x"66686B6E", x"6F6F6E6E", x"6F707173", x"76777674", x"78787A7E", x"82848382",
									 -- x"85848587", x"8887898B", x"8A8A8C8F", x"908F9195", x"9095999C", x"A0A0A2A9", x"A3A6A7A8", x"ABA8A8AE",
									 -- x"ADACAEB3", x"B5B2B1B4", x"B8B2AEAF", x"AEABACAF", x"ADA8A6A7", x"A8A5A4A5", x"A9A7A6A7", x"A6A2A0A0",
									 -- x"9D9A999B", x"9A969596", x"94929192", x"918D8C8D", x"88898A8B", x"8A898988", x"86837F7D", x"7C7B7D7F",
									 -- x"7D7F7E79", x"7371706F", x"71737372", x"72747471", x"76716E70", x"72716E6E", x"6B70726F", x"6F73716A",
									 -- x"7072767C", x"7F808284", x"898B8C8A", x"888B9196", x"979B9FA1", x"A4A8A9A9", x"AEB7BDBF", x"C1BFC0C5",
									 -- x"C8CCD0D3", x"D5D8DDE1", x"E7ECEEEA", x"E6E6E9EB", x"ECEBE9E6", x"E3E2E0DD", x"E0E0E2E7", x"EDF1F0EE",
									 -- x"EFEDEAE7", x"E3E2E3E5", x"E7E6E6E6", x"E5E3E0DE", x"DAD9D4CF", x"CDCECECB", x"C8CACAC6", x"C2C2C1BF",
									 -- x"C5C0BBB8", x"B7B6B4B2", x"B4B6B5B5", x"B6B3B3B7", x"B8BAB9B8", x"B8B5B6BC", x"C4C2BEBE", x"BFBAB7BB",
									 -- x"C0C4C1B7", x"B3B5B2AB", x"A8A7A5A1", x"9C9A9B9D", x"9A9A9292", x"94959995", x"97999DA2", x"A3A3A3A4",
									 -- x"A7AAB0B6", x"BEC3C1BD", x"C1BEBBBA", x"BBBDBDBC", x"C4C8CED4", x"D8DADBDC", x"D6D4D3D4", x"D4D1CFCF",
									 -- x"C7C7C5BE", x"B7B1B0B1", x"ACA6A4A8", x"A7A0A0A6", x"ABA8A7A9", x"AAA9A9AB", x"A8AAADAA", x"A5A8AAA6",
									 -- x"A5A6A5A2", x"A1A3A4A3", x"A7A39D99", x"95918F90", x"8D868687", x"827D7D7C", x"7A797979", x"79787877",
									 -- x"78757372", x"716E6D6E", x"6F6F6967", x"69696667", x"615F5D5E", x"60605C59", x"58535154", x"55525051",
									 -- x"4D4B4948", x"4B4E4E4B", x"46454443", x"42413E3B", x"41403F3E", x"3C3A3837", x"34343434", x"3432302F",
									 -- x"2D2E2D2B", x"2B2B2825", x"27262524", x"23232425", x"21212223", x"201D1D1F", x"24232221", x"22232322",
									 -- x"E5E7E7E7", x"E8EAE9E6", x"E5E5E6E6", x"E6E6E6E5", x"E4E5E6E6", x"E6E6E6E5", x"E4E4E4E3", x"E3E2E1E1",
									 -- x"E2E3E3E4", x"E4E3E1E0", x"DEDEDCD9", x"D6D5D7D9", x"D1D3D3D2", x"CFCCC9C7", x"C7C7C6C3", x"C3C5C4C1",
									 -- x"BFBCB5AE", x"A8A39D99", x"95908B8B", x"8A868281", x"7C7C7976", x"75767572", x"70706F70", x"7273726F",
									 -- x"70717272", x"72737475", x"7473706E", x"6C6A6968", x"69696868", x"67666564", x"68686866", x"64636466",
									 -- x"66646364", x"66656667", x"6664686A", x"68676969", x"696D7275", x"75747272", x"75777A7D", x"7F808284",
									 -- x"85858687", x"8785878A", x"8B8A8C91", x"8F8B8C91", x"9292959B", x"9E9E9EA0", x"A3A3A3A4", x"A5A7A9AA",
									 -- x"ABAAABAD", x"B0B2B1B1", x"B1B3B1AC", x"A9A9AAAA", x"A9A8A6A5", x"A4A4A5A5", x"A6A3A2A0", x"9E9F9E99",
									 -- x"97999893", x"90919394", x"958F8C8D", x"8F8F8C8A", x"8A8B8A88", x"88888786", x"8584817D", x"7B7C7C7B",
									 -- x"79787775", x"75777674", x"72737475", x"75757576", x"76757777", x"75727173", x"70727474", x"72717274",
									 -- x"747A7E7D", x"7E858C8E", x"8E909394", x"9597999C", x"A1A1A4A9", x"ACAEB2B6", x"B9BFC4C5", x"C5C8CACB",
									 -- x"D3D6D9DB", x"DCDFE4E8", x"EFF3F5F1", x"EDECEDED", x"F2F0EEEA", x"E7E4E2E1", x"E3E4E5E9", x"EFF2F0EC",
									 -- x"EFECE9E6", x"E5E5E6E6", x"E6E7E7E6", x"E6E5E2DF", x"DBDAD6D1", x"CFD0CFCD", x"CFCDCDCE", x"CDCCCBCC",
									 -- x"CBCAC8C4", x"C1BFBDBB", x"B9BBBCBB", x"BABBBCBB", x"BAB7BABE", x"BAB8BBBF", x"C4C2C4C8", x"C3BAB9C0",
									 -- x"BDC1C3C2", x"BFB9B2AC", x"A8AAA7A0", x"9C9B9895", x"97959494", x"92919294", x"9396999C", x"9EA0A2A4",
									 -- x"A3A6ACB5", x"BABBBABA", x"BBBDBDBB", x"BBBCBEBE", x"C2C5CBD3", x"D8D8D6D6", x"D2CFCECE", x"CECCCBCB",
									 -- x"CBC6C1BD", x"B8B2ADAB", x"A8A5A4A5", x"A5A3A3A5", x"A0A9ABA7", x"A6A7A7A9", x"AAACACA8", x"A5A5A6A6",
									 -- x"A1A3A5A5", x"A3A5A9AF", x"ADABA49D", x"9B9A958D", x"8C837D7F", x"827F7976", x"79777576", x"77767473",
									 -- x"6E70706D", x"6C6D6D6C", x"686A6B68", x"66666665", x"5F60615E", x"5B5A5A5B", x"5B555555", x"514E5052",
									 -- x"4D4D4D4C", x"4E504D49", x"46474643", x"4343413E", x"41403F3E", x"3D3C3A39", x"38383837", x"35333332",
									 -- x"2B2F2F2C", x"2B2C2B27", x"29272628", x"28252425", x"24212021", x"21202022", x"22212122", x"25262523",
									 -- x"E6E6E6E5", x"E5E7E7E5", x"E6E6E6E6", x"E6E6E6E5", x"E6E6E7E7", x"E7E6E6E5", x"E4E4E3E3", x"E2E2E1E1",
									 -- x"E0E0E1E2", x"E2E2E1DF", x"DCDBDAD8", x"D6D5D5D6", x"D5D5D4D1", x"CECBC9C8", x"C4C6C6C4", x"C3C3C3C1",
									 -- x"BBB9B4AE", x"A9A5A09B", x"97928D8B", x"8985817E", x"7E7C7774", x"74757370", x"6F6F6F70", x"706F6F6E",
									 -- x"70707171", x"70707172", x"72706C6B", x"6B6A6865", x"64646465", x"66676766", x"62636363", x"62616162",
									 -- x"62606061", x"62616162", x"62606468", x"66676B6B", x"6B6C6E6F", x"6F707172", x"7274777A", x"7C7D7F81",
									 -- x"85858687", x"8685878A", x"89888A8E", x"8F8D8D8F", x"93929497", x"99999A9C", x"9F9FA0A1", x"A3A5A7A9",
									 -- x"AAAAAAAA", x"AAABACAD", x"AEB0B0AC", x"A9A9A9A9", x"A6A6A6A5", x"A5A3A2A1", x"A3A1A1A0", x"9D9E9D97",
									 -- x"9595938F", x"8E90908E", x"908B888A", x"8C8B8988", x"87878787", x"898A8885", x"8384827E", x"7C7B7A77",
									 -- x"79797876", x"77777674", x"76777879", x"7A7A7978", x"7979797B", x"7A777779", x"75757676", x"7677797A",
									 -- x"767E8586", x"898F9495", x"98999B9C", x"9C9DA1A3", x"A9AAACB1", x"B4B5B8BC", x"BEC1C4C7", x"CBCFD2D2",
									 -- x"DADCE0E2", x"E3E6EBEF", x"F4F7F9F6", x"F3F2F2F1", x"F4F3F0ED", x"EBE9E7E7", x"E7E8E9EB", x"EFF1EFEB",
									 -- x"ECEBEAE9", x"E8E7E5E4", x"E8EAEBEB", x"EAE9E5E1", x"DDDCD9D5", x"D4D5D5D3", x"D3D2D3D4", x"D4D2D1D2",
									 -- x"CECECDCB", x"C8C6C4C3", x"BDBFC0BF", x"BFC1C2C1", x"BBB7B9BC", x"B9B8BEC2", x"C5C2C3C5", x"C2BBB8BB",
									 -- x"B8BEC4C3", x"BDB6AFAA", x"A8A7A49E", x"9A979491", x"8F8F9092", x"92919192", x"97989999", x"9899999A",
									 -- x"A0A3A9B0", x"B3B4B6B9", x"BABBBAB8", x"B7BABCBD", x"C2C3C7CD", x"D1D1D0D0", x"D3D1CFCC", x"C8C5C6C8",
									 -- x"C9C4BEBA", x"B6B1ADAC", x"A6A4A2A2", x"A19FA0A1", x"9FA7A9A6", x"A7A9A9AB", x"A8A9A9A8", x"A8A8A8A6",
									 -- x"A0A5ADB2", x"B2B1B0B0", x"ACA9A39E", x"9D9D958C", x"8A848284", x"837D7775", x"79777474", x"73727170",
									 -- x"6A6C6B6A", x"696B6C6B", x"686A6A67", x"65666665", x"5C5C5D5B", x"59585859", x"57514F52", x"5353524D",
									 -- x"50504E4D", x"4F514F4B", x"494A4947", x"47484745", x"4141403F", x"3E3D3C3A", x"3A3A3937", x"35353535",
									 -- x"2C2E2D2A", x"2B2E2C28", x"29272729", x"29262526", x"26252627", x"25232224", x"22212224", x"27292928",
									 -- x"E4E6E6E5", x"E5E6E4E2", x"E5E5E5E5", x"E5E5E4E4", x"E6E6E6E6", x"E6E5E5E5", x"E4E4E3E2", x"E2E1E1E1",
									 -- x"DEDEDFE0", x"E1E1E1E0", x"DAD9D8D8", x"D7D6D5D4", x"D6D3D0CC", x"C9C6C5C5", x"C1C3C4C3", x"C2C1C0BF",
									 -- x"B9B7B3AE", x"AAA7A29D", x"99948F8C", x"8A85807E", x"7E7A7571", x"7172706D", x"6E6D6E70", x"6F6C6D70",
									 -- x"6F6F6F6F", x"6E6D6E6E", x"706D6968", x"69696663", x"64636363", x"64646362", x"5E5E5F61", x"61615F5E",
									 -- x"605E5E5F", x"5F5E5E5E", x"605E6165", x"64656969", x"696A6B6B", x"6A6C6E70", x"6F727577", x"797B7C7D",
									 -- x"7E7F8082", x"82818386", x"8888888A", x"8C8D8C8B", x"91919293", x"93939598", x"9A9B9C9E", x"A0A3A5A7",
									 -- x"A8A9A9A7", x"A5A6A8AB", x"AAADADAB", x"A9A8A8A8", x"A6A6A5A4", x"A4A2A09E", x"A09FA1A0", x"9B9B9A95",
									 -- x"9794918F", x"90918F8B", x"8B888688", x"88878686", x"86868586", x"898B8884", x"81838381", x"7F7D7A77",
									 -- x"7B7C7B79", x"797A7876", x"7A7B7D7F", x"80807F7E", x"7F7E7D7E", x"7F7D7D7D", x"7B7A7A7B", x"7D7F8181",
									 -- x"83888B8A", x"8C939A9D", x"A1A2A3A3", x"A2A4A8AC", x"B0B1B5B9", x"BCBDC0C2", x"C4C4C5C9", x"D0D6D9D8",
									 -- x"DEE1E5E7", x"E9ECF1F4", x"F6F9FBFB", x"FBFAF8F6", x"F6F4F1F0", x"EFEEEEED", x"EBEDEDED", x"EEEFEDEA",
									 -- x"EEEDECEA", x"E9E7E5E4", x"E7E9EBEC", x"EBEAE6E1", x"DEDDDBD8", x"D7D8D8D7", x"D7D7D7D9", x"D8D6D4D4",
									 -- x"D3D3D3D2", x"D0CECCCB", x"C4C5C5C3", x"C3C5C5C4", x"BDBABCBE", x"BABABEC0", x"BEBEC0C2", x"C2BFBBBA",
									 -- x"B5BDC3C2", x"BBB4AFAD", x"A8A4A09C", x"9893908F", x"918F8F90", x"908E8D8D", x"91929394", x"9597999B",
									 -- x"9FA2A7AB", x"ADAFB3B8", x"B4B5B4B3", x"B5BBC0C2", x"C5C4C6C9", x"CCCCCCCD", x"D2D1CEC9", x"C2BDC0C5",
									 -- x"C5C0B9B5", x"B1ADABAB", x"A4A3A2A0", x"9E9C9D9F", x"9FA5A6A4", x"A7A8A8AA", x"A6A6A7A8", x"AAABA8A5",
									 -- x"A5A9AEB2", x"B4B4B3B3", x"ACAAA6A2", x"A2A0978D", x"88878687", x"847E7B7B", x"78767370", x"6E6D6C6B",
									 -- x"6B6B6967", x"66676767", x"67686765", x"63646464", x"5B5C5C5C", x"5B595756", x"57535253", x"54575750",
									 -- x"5452504F", x"5152514E", x"4D4D4C4B", x"4B4C4C4A", x"44444343", x"4241403E", x"3C3A3835", x"34343535",
									 -- x"2F302E2B", x"2C2F2D2A", x"29282829", x"28262525", x"25262829", x"29262425", x"27262526", x"28292928",
									 -- x"E2E4E6E7", x"E7E7E3E0", x"E3E3E3E3", x"E3E2E2E2", x"E4E4E4E4", x"E4E4E4E4", x"E4E4E3E2", x"E2E2E2E2",
									 -- x"DEDEDEDF", x"E0E1E1E0", x"DCDAD8D8", x"D7D6D4D3", x"D2CFCAC7", x"C4C1C0C1", x"C0C0C0C0", x"C0BFBCB9",
									 -- x"B8B6B2AD", x"A9A6A29E", x"99958F8C", x"8A86827E", x"7B797571", x"6F6F6E6C", x"6C6A6B6E", x"6E6C6C70",
									 -- x"6E6E6E6D", x"6C6B6C6D", x"6E6C6967", x"67666463", x"64646362", x"61605F5E", x"5E5E5F60", x"62615F5D",
									 -- x"5F5D5C5D", x"5D5C5C5D", x"625F6164", x"62626564", x"6466696A", x"6A6A6A6B", x"6C6F7273", x"75777878",
									 -- x"76787A7B", x"7C7D8082", x"86888988", x"898A8A87", x"8D8E8F90", x"8F8F9295", x"93959799", x"9B9EA1A3",
									 -- x"A6A6A6A5", x"A5A5A7A8", x"A8A9AAAA", x"A9A8A8A8", x"ABA9A5A3", x"A2A1A09F", x"9D9D9F9D", x"99989894",
									 -- x"97949190", x"9292908C", x"8A888788", x"88868687", x"88888786", x"88898784", x"81828483", x"82807E7B",
									 -- x"7F7F7E7C", x"7B7C7D7B", x"7B7E8184", x"85858686", x"85838181", x"82828180", x"807F7E80", x"83868686",
									 -- x"8C8E8F8E", x"90979EA2", x"A6A7A8A8", x"A8ABB0B4", x"B7B9BDC1", x"C4C5C7C9", x"CCCBCBCE", x"D5DBDEDE",
									 -- x"E1E4E9EC", x"EFF1F4F6", x"F5F6F9FC", x"FFFFFDFA", x"F6F4F1F0", x"F1F2F2F2", x"F1F3F2F0", x"EFF0F0EF",
									 -- x"F5F1EDE9", x"E7E7E7E7", x"E4E7E9EA", x"EAE9E6E1", x"DFDEDCDA", x"DADAD9D8", x"DBDADBDC", x"DBD7D5D4",
									 -- x"D7D6D6D6", x"D5D2CFCF", x"CCCDCBC9", x"C7C7C5C2", x"BEBCBFC1", x"BCB8B9B8", x"B7BBBFC1", x"C1C0BDBA",
									 -- x"B5BABEBB", x"B6B2B0AF", x"A7A19C9B", x"98928F8F", x"95928F8E", x"8D8C8C8D", x"94949494", x"94949494",
									 -- x"9C9EA3A7", x"AAABAFB3", x"B1B2B1B1", x"B5BDC3C6", x"C7C6C6C8", x"CACACBCC", x"CECCC9C5", x"BEBBBDC2",
									 -- x"C1BCB5B1", x"ADA9A6A6", x"A2A2A2A0", x"9D9C9EA0", x"9FA4A4A3", x"A6A6A4A4", x"A5A5A5A7", x"A8A9A7A5",
									 -- x"AAABADAE", x"AFB1B0AF", x"AAABABAA", x"A8A49A91", x"8E8C8A88", x"84807F81", x"7A7A7772", x"6F6E6C6B",
									 -- x"6D6B6866", x"65666666", x"65656463", x"62636363", x"61606061", x"605C5856", x"59595A56", x"52565A58",
									 -- x"55545352", x"53535250", x"50504F4E", x"4D4C4B49", x"46454545", x"45434240", x"3D3B3936", x"35343434",
									 -- x"3233322F", x"2F2F2E2B", x"2C2C2C2B", x"29272626", x"25252629", x"2B2A2826", x"2A292828", x"292A2929",
									 -- x"DFE1E3E3", x"E4E4E2E0", x"E1E1E1E1", x"E1E1E1E0", x"E2E2E2E2", x"E3E3E3E4", x"E4E4E3E3", x"E2E2E1E1",
									 -- x"DEDDDDDD", x"DEDFDFDE", x"DDDBD8D7", x"D6D5D3D1", x"CECAC7C6", x"C3C0BEBE", x"BFBCBABB", x"BCBBB7B3",
									 -- x"B5B3AFAA", x"A7A5A19E", x"97938E8B", x"8886817D", x"76787672", x"6F6E6D6C", x"6D69686B", x"6D6B6A6B",
									 -- x"6B6B6A69", x"69696A6B", x"6B6B6966", x"64626262", x"60606060", x"6161605F", x"605F5F5F", x"60615F5E",
									 -- x"5D5B5959", x"5A5A5B5C", x"615E6062", x"61616261", x"61646768", x"68686868", x"696C6F6F", x"6F727372",
									 -- x"73757778", x"797B7D7F", x"83868988", x"87888989", x"898C8E8E", x"8D8D8F91", x"8C8E9193", x"94979A9C",
									 -- x"A2A2A2A3", x"A4A5A4A3", x"A6A6A7A7", x"A7A7A8A9", x"ABA9A5A3", x"A2A19F9E", x"9D9C9D9B", x"96969793",
									 -- x"92919090", x"908F8E8D", x"8A898989", x"88868587", x"87888886", x"84858685", x"83848485", x"8482807F",
									 -- x"8282807D", x"7D7F8181", x"7D828789", x"88888A8C", x"8A898787", x"87888785", x"86848486", x"898B8A88",
									 -- x"8A8F9598", x"9B9FA3A4", x"A9ABACAE", x"AFB4BABE", x"C2C5C9CC", x"CECFCFCF", x"D2D1D2D5", x"D9DEE2E4",
									 -- x"E6EAEFF3", x"F5F7F8F9", x"F5F5F6FB", x"FFFFFDFB", x"F6F4F2F2", x"F4F6F6F6", x"F7F8F7F4", x"F2F4F6F6",
									 -- x"F8F3EDE8", x"E6E6E7E8", x"E4E6E8E8", x"E9E9E7E4", x"E0DFDEDE", x"DEDDDCDC", x"DEDDDEDF", x"DEDAD8D8",
									 -- x"D7D6D6D8", x"D7D4D2D2", x"D3D3D2CF", x"CCCAC6C2", x"BFBDBFC0", x"BAB6B5B3", x"B5BBC0C0", x"BFBDBAB6",
									 -- x"B5B7B7B5", x"B2B0AEAB", x"A69F9A99", x"97928E8E", x"928F8D8D", x"8E8E8F90", x"90919192", x"93939393",
									 -- x"97989CA2", x"A6A8A9AB", x"B2B3B2B3", x"B7BEC3C5", x"C5C4C4C7", x"C9C8C8C9", x"C6C4C2C0", x"BEBCBDC0",
									 -- x"BEB9B4B0", x"ABA6A2A0", x"9FA0A09D", x"9B9C9FA1", x"9FA3A3A3", x"A5A4A0A0", x"A2A2A3A4", x"A4A5A5A6",
									 -- x"A7ABAFB1", x"B2B1ABA5", x"A3A8ADAE", x"ABA49C96", x"95928E8B", x"86828080", x"7F81807B", x"76757371",
									 -- x"6E6B6867", x"67686A6B", x"66666667", x"67676667", x"68656363", x"615D5B5B", x"595A5C58", x"53575B58",
									 -- x"56555556", x"56555352", x"52515151", x"504D4B49", x"47474646", x"45444240", x"413F3D3B", x"3A383635",
									 -- x"31333433", x"312F2E2C", x"2E2F2F2D", x"2C2B2B2A", x"2A282729", x"2D2E2B27", x"2A2A2A2B", x"2C2E2E2F",
									 -- x"DDDDDCDA", x"DCDFE0DF", x"DEDFDFE0", x"E0E0E0E0", x"E0E0E0E0", x"E1E2E2E3", x"E2E2E2E2", x"E2E1E0E0",
									 -- x"DDDCDBDA", x"DBDCDCDC", x"DBDAD8D6", x"D5D3D1D0", x"CBC6C4C4", x"C2BEBABA", x"BCB8B5B6", x"B7B5B1AE",
									 -- x"B0AEABA6", x"A4A3A09D", x"95928D89", x"8785807C", x"73757471", x"6E6D6C6A", x"6F6C6969", x"6A6A6866",
									 -- x"68686766", x"66666869", x"68696865", x"615F5F60", x"5F5E5E5F", x"60605F5E", x"605F5E5E", x"5E5E5D5D",
									 -- x"5E5B5959", x"59595B5C", x"5B585B5F", x"5F606261", x"60626363", x"63646668", x"6A6D6E6C", x"6C6F706E",
									 -- x"71737574", x"74767879", x"7D818486", x"8686888B", x"888A8C8B", x"8B8B8B8A", x"898B8E90", x"90929597",
									 -- x"9B9B9C9E", x"A0A09E9B", x"A3A2A2A4", x"A5A5A6A7", x"A6A5A4A5", x"A4A29D9A", x"9D9B9B99", x"95969692",
									 -- x"908F8F8F", x"8E8D8D8E", x"8A898889", x"88868586", x"85878784", x"83848687", x"87868586", x"85838182",
									 -- x"83838280", x"80838687", x"85898E8F", x"8D8D8E91", x"8F90908F", x"9091918F", x"8D8C8B8D", x"8F908F8D",
									 -- x"9194989B", x"9EA2A6A8", x"ACAEB1B4", x"B7BCC2C6", x"CCD0D4D5", x"D6D6D5D4", x"D3D4D6D9", x"DCDFE4E8",
									 -- x"EBEEF2F6", x"F8F9F9FA", x"F8F6F6FA", x"FEFEFDFB", x"F9F7F5F6", x"F8FAFAF9", x"F8F9F7F5", x"F4F6F8F8",
									 -- x"F6F3EFEB", x"E8E7E7E7", x"E5E7E7E7", x"E7E8E7E4", x"E0DFDFE0", x"E1DFDEDE", x"DEDDDDDE", x"DDDBDADA",
									 -- x"D7D5D6D8", x"D8D5D5D6", x"D4D4D2CF", x"CECCC8C3", x"C5C2C2C0", x"BAB9B9B7", x"B2B7BBBB", x"BAB9B8B7",
									 -- x"B6B6B5B4", x"B3B1ABA6", x"A59F9996", x"95938F8C", x"8F8E8E90", x"918F8D8C", x"88888A8C", x"90939495",
									 -- x"9494989E", x"A3A5A6A7", x"ACAEB0B3", x"B9BFC3C4", x"C2C1C2C5", x"C6C5C4C5", x"BDBBBABB", x"BCBCBCBC",
									 -- x"BBB6B2AE", x"AAA49F9D", x"9B9C9C99", x"989A9D9E", x"9FA3A2A2", x"A4A29FA0", x"9F9E9FA0", x"A1A1A3A6",
									 -- x"A3A9AEAF", x"B0AFA9A3", x"9DA3AAAC", x"A9A29C99", x"9291908F", x"8D8A8785", x"85888882", x"7D7B7A78",
									 -- x"77726D6B", x"6B6B6C6D", x"6D6C6D70", x"706F6D6D", x"6C676361", x"5F5D5F63", x"5C5A5B5D", x"5D5E5D57",
									 -- x"5857585A", x"5A585656", x"55545455", x"54514F4E", x"4C4C4B4B", x"49474442", x"42413F3E", x"3D3B3735",
									 -- x"30323434", x"3332302E", x"2D2E2E2C", x"2A2B2C2D", x"2F2B2828", x"2B2E2B26", x"2E2E2E2E", x"2F303232",
									 -- x"D8D9D7D6", x"D8DBDCDB", x"DBDBDCDD", x"DDDEDEDE", x"DEDEDDDD", x"DEDEDFE0", x"E0E0E1E1", x"E1DFDEDD",
									 -- x"DCDBD9D9", x"DADADBDB", x"D9DAD9D8", x"D5D3D1D0", x"CBC6C3C4", x"C2BCB8B7", x"B7B4B2B2", x"B0AEADAE",
									 -- x"ABABA8A5", x"A2A09C98", x"94928D89", x"8887837E", x"78777472", x"71716F6C", x"70716F6A", x"6A6B6A66",
									 -- x"68676766", x"65666769", x"68676664", x"61605F60", x"5F5F5E5E", x"5E5D5C5B", x"5D5D5D5C", x"5B5B5B5B",
									 -- x"5D5B5A5A", x"5B59595A", x"5553575C", x"5D5E5F5D", x"5E5E5F5F", x"5F616467", x"696C6C69", x"686B6C6A",
									 -- x"6B6E706F", x"6F727474", x"78787B80", x"82818386", x"86888988", x"87888886", x"86898C8D", x"8C8D8F91",
									 -- x"92939698", x"9A9A9998", x"9E9D9EA1", x"A2A2A2A3", x"A3A2A2A4", x"A5A39E9A", x"9D9A9A99", x"96969690",
									 -- x"918F8E8F", x"8E8C8C8E", x"8A888889", x"89888686", x"86878785", x"85878888", x"89878788", x"87858485",
									 -- x"84868685", x"86898C8D", x"90919394", x"95959596", x"95989998", x"98999998", x"95949494", x"96979696",
									 -- x"9D9D9C9D", x"A0A4AAAF", x"B2B5B9BC", x"C0C4C9CD", x"D2D6DADC", x"DCDDDBD9", x"D8D8DBDF", x"E1E3E7EB",
									 -- x"F0F1F3F6", x"F7F9FAFA", x"FBF7F6F8", x"FBFCFCFD", x"FDFAF8F9", x"FBFDFCFB", x"F8F8F8F6", x"F6F7F7F6",
									 -- x"F7F4F1EE", x"EDEBEAEA", x"E9EAEAE9", x"E9E9E7E4", x"E4E2E2E4", x"E3E0DEDE", x"DEDCDBDB", x"DAD8D7D8",
									 -- x"D7D5D5D8", x"D8D5D5D8", x"D3D2D0CD", x"CCCCC9C6", x"CAC6C6C3", x"BEBDBEBB", x"B1B1B2B3", x"B4B4B5B6",
									 -- x"B4B3B2B0", x"AFAEA9A4", x"A29E9895", x"9697948F", x"94929192", x"918D8987", x"8C8A8887", x"898B8C8C",
									 -- x"9393969B", x"9FA1A5A8", x"A7AAAEB2", x"B8BDBEBD", x"BEBCBDBF", x"BFBEBCBD", x"B7B5B5B6", x"B8B7B6B7",
									 -- x"B5B1ADAA", x"A7A29E9C", x"9A9A9996", x"95989A9A", x"9FA2A09E", x"A09E9DA0", x"9E9B9A9D", x"9F9FA0A1",
									 -- x"A2A6A9A8", x"A8AAA8A4", x"9DA1A6A8", x"A49F9A98", x"91929393", x"9291908F", x"8D909089", x"83828180",
									 -- x"807A7472", x"72717274", x"74747679", x"7A777372", x"6F6A6765", x"625F6166", x"605D5F64", x"6362615D",
									 -- x"5C5B5B5D", x"5D5C5B5C", x"5B595859", x"58565455", x"5151504F", x"4D4A4644", x"43413F3E", x"3E3C3937",
									 -- x"34333335", x"37363330", x"2E302F2B", x"292A2C2D", x"2F2E2B29", x"2A2C2B28", x"32313131", x"31313233",
									 -- x"D4D6D7D7", x"D8DAD9D7", x"D7D8D9DA", x"DADBDBDB", x"DBDBDBDA", x"DADBDBDC", x"DEDFE0E0", x"E0DEDCDB",
									 -- x"DCDBDAD9", x"DADBDCDC", x"D8DADBDA", x"D7D4D2D1", x"D0CAC6C6", x"C4BDB8B8", x"B3B2B1AF", x"ACA9AAAE",
									 -- x"AAAAA8A5", x"A29E9893", x"93918E8A", x"8A8B8883", x"817E7976", x"78797671", x"7175746D", x"6B6E6E6A",
									 -- x"69696867", x"66676869", x"69676564", x"63626160", x"5D5D5C5D", x"5D5D5C5B", x"5A5C5D5C", x"5B595A5B",
									 -- x"5A595859", x"59575656", x"5451555A", x"5A5A5B58", x"5A5B5C5D", x"5E5F6264", x"65686763", x"63666765",
									 -- x"676B6D6C", x"6D717474", x"7471737A", x"7E7C7C80", x"84868584", x"85878684", x"82858788", x"8786888B",
									 -- x"8B8E9294", x"95969798", x"9A999B9F", x"A09F9E9F", x"A3A1A1A2", x"A4A4A19E", x"9C9A9A99", x"9797958F",
									 -- x"918E8C8D", x"8D8B8B8C", x"8A88888A", x"8B898887", x"89898988", x"898A8987", x"8988888B", x"8B888889",
									 -- x"86898B8B", x"8C8F9192", x"96959698", x"9B9D9C9A", x"9A9E9F9D", x"9C9D9D9B", x"9B9A9999", x"9A9B9C9C",
									 -- x"9E9FA2A6", x"A9ADB1B4", x"B9BDC1C5", x"C8CCD1D4", x"D4DADEE0", x"E1E2E1DE", x"DFDFE1E5", x"E8E9EBEE",
									 -- x"F5F5F5F6", x"F7F9FBFD", x"FBF7F5F7", x"FAFBFDFF", x"FEFCFAFB", x"FDFEFDFB", x"FAFBFBFA", x"FAFBF9F6",
									 -- x"FAF7F3F0", x"EFEFEFF0", x"EEEFEFEE", x"EEEDEAE7", x"EBE9E8E9", x"E7E3DFDF", x"E1DEDCDA", x"D8D6D5D7",
									 -- x"D9D6D5D8", x"D7D4D4D7", x"D5D3D0CD", x"CDCECCC9", x"C9C7C7C5", x"C0BEBCB8", x"B6B0ACAE", x"AFAFB0B2",
									 -- x"AFAEABA8", x"A8A8A7A4", x"A09D9895", x"989C9994", x"99959291", x"908D8988", x"88858383", x"868A8D8F",
									 -- x"90909396", x"989CA2A9", x"A8ABAEB2", x"B5B7B5B2", x"B8B6B6B7", x"B7B5B3B4", x"B5B3B2B3", x"B3B2B2B2",
									 -- x"B0ACA8A6", x"A39F9C9B", x"9B9A9794", x"94979897", x"A0A19E9B", x"9B99999E", x"9F9B989B", x"9E9E9D9C",
									 -- x"9EA4A8A7", x"A7A8A6A2", x"A2A3A5A5", x"A19C9896", x"99999996", x"93929496", x"9599978F", x"89898988",
									 -- x"827C7777", x"787A7C7F", x"79787B7F", x"7F7B7674", x"706E6E6D", x"69626165", x"62606467", x"625F6264",
									 -- x"605E5D5F", x"5F5E5E60", x"605D5A5B", x"5A585759", x"5251504E", x"4C484542", x"45434140", x"41403D3B",
									 -- x"3B363335", x"3A3A3631", x"3435332E", x"2B2C2E2F", x"3031302D", x"2C2D2E2D", x"2F2F3030", x"31333537",
									 -- x"CED0D3D4", x"D5D6D7D8", x"D3D4D5D6", x"D5D6D8DA", x"D9DAD9D6", x"D7DBDCDB", x"DFDFDFDF", x"DEDEDCDB",
									 -- x"DBDAD9D8", x"D7D7D8DB", x"DADADAD9", x"D7D6D4D3", x"D1CFCCC9", x"C4C0BCBA", x"B9B1ADB0", x"B0ABA9AC",
									 -- x"AAA5A4A3", x"9E9B9994", x"93919090", x"8E8C8B8C", x"89878380", x"7F7F7D7A", x"78777778", x"7672706F",
									 -- x"6B696664", x"666A6B69", x"6A6A6966", x"63626263", x"605F5C5A", x"5B5C5D5D", x"5C5C5D5C", x"5C5C5C5D",
									 -- x"5A585758", x"59595653", x"57555455", x"595B5A58", x"54585B59", x"5A5E5F5E", x"60626462", x"605F6163",
									 -- x"65676867", x"6B71726F", x"73706F72", x"76787A7B", x"787A7F7D", x"80878381", x"83828182", x"85878887",
									 -- x"8A8A8C8E", x"9090908F", x"9092979B", x"9B989A9E", x"9EA0A3A4", x"A2A09E9E", x"9A999896", x"95949393",
									 -- x"8F8E8E8F", x"8E8C8B8B", x"8B8A8B8C", x"8B8A8B8E", x"8D8A8A8D", x"8D8A898C", x"8E8D8C8B", x"8B8C8E8F",
									 -- x"918E8D90", x"93959799", x"989A9C9D", x"9FA1A3A4", x"A5A3A3A6", x"A8A7A5A4", x"A3A09F9F", x"A0A0A2A5",
									 -- x"A2A6ABAD", x"AFB2B9BE", x"C0C2C6CA", x"CBCDD2D9", x"DBE0E2E2", x"E3E6E6E4", x"E4E3E2E4", x"E8EDF1F3",
									 -- x"F6F5F4F4", x"F6F8F9FA", x"F9F9F9FA", x"FCFEFEFF", x"FDFDFCFC", x"FDFEFEFE", x"FDFCFCFD", x"FDFDFBF9",
									 -- x"FBF8F5F3", x"F4F4F4F3", x"F1F4F5F2", x"EFEFEFEF", x"EFEDEBEA", x"E8E6E3E1", x"E0DEDBD8", x"D6D6D5D5",
									 -- x"D5D5D7D9", x"D9D6D4D4", x"CED2D2CC", x"C8C9CCCF", x"CCC8C8C9", x"C4BEBBB7", x"B3AFABA9", x"ABADAEAE",
									 -- x"AAA8A6A3", x"A09F9FA1", x"9E9C9A98", x"97989796", x"9594918D", x"8B89847E", x"85828182", x"8383868A",
									 -- x"8890928F", x"92979A9E", x"A3A6ABB1", x"B4B3B1AF", x"B2B5B2B4", x"B2AEB2B0", x"B1B1AFAF", x"B0B2B0AD",
									 -- x"ADAAA8A7", x"A59F9895", x"93959694", x"8F8C9096", x"969B9D9B", x"9A9B9996", x"9C9B9A97", x"9696999B",
									 -- x"9DA5A5A3", x"A7A8A6A9", x"A5A1A0A4", x"A49D9693", x"99999A98", x"94919396", x"9A949697", x"8F8F8F87",
									 -- x"8E8E8A86", x"84868685", x"81828886", x"827F7776", x"74716D6A", x"6B6D6B66", x"68696A6A", x"6A6A6867",
									 -- x"64626265", x"64615F5F", x"63605D5D", x"5E5E5B59", x"5A56524F", x"4E4E4C4A", x"49494743", x"4242423F",
									 -- x"3C3B3937", x"38393733", x"36333233", x"33302D2D", x"2F313231", x"30313130", x"31333536", x"35343536",
									 -- x"CCCED0D1", x"D1D1D2D2", x"D0D1D2D3", x"D3D4D6D7", x"D5D5D5D4", x"D4D6D7D7", x"DBDBDBDC", x"DCDCDBDA",
									 -- x"D9D8D7D5", x"D5D6D7D8", x"D8D8D8D8", x"D7D6D5D4", x"D1D1CFCC", x"C7C2BFBC", x"B9B4B0B0", x"AFABAAAC",
									 -- x"A9A4A4A2", x"9E9C9A95", x"95929190", x"8F8D8D8E", x"8B898785", x"83817F7E", x"7A787777", x"76737070",
									 -- x"6F6E6D6B", x"6B6D6D6B", x"6C6C6B69", x"67656464", x"615F5D5B", x"5B5B5C5B", x"595A5B5B", x"5B5B5B5B",
									 -- x"58585858", x"58575655", x"53535354", x"55565555", x"53565858", x"58595A5A", x"5D5F6060", x"5F5F6062",
									 -- x"60656868", x"6B6D6C68", x"6C6A696C", x"6F727476", x"78787B77", x"787E7A79", x"7F7E7E80", x"83858585",
									 -- x"87878889", x"8B8C8D8D", x"91919294", x"9596989B", x"9B9C9D9F", x"A09F9D9C", x"9A999896", x"9492908F",
									 -- x"908E8E8F", x"8F8D8D8E", x"8D8D8E90", x"8F8E8D8F", x"8F8D8D90", x"918F8F92", x"91919090", x"90919192",
									 -- x"92919296", x"999A9C9E", x"9D9FA0A2", x"A4A6A9AB", x"ACA9A8AB", x"ACABA9A8", x"A7A5A4A5", x"A5A5A7A9",
									 -- x"ABADB0B3", x"B6BABEC1", x"C5C7CBCE", x"D0D1D7DD", x"DCE1E3E3", x"E4E8E8E6", x"E7E6E4E4", x"E7ECF0F2",
									 -- x"F3F2F2F3", x"F5F8F9FA", x"F8F9FAFC", x"FDFEFEFE", x"FDFCFCFC", x"FDFEFEFE", x"FEFDFCFC", x"FDFDFCFB",
									 -- x"FCF9F7F6", x"F6F7F6F5", x"F4F6F5F2", x"EFEFEEED", x"EEEDECEB", x"EAE8E5E2", x"DFDDD9D7", x"D6D6D5D5",
									 -- x"D5D6D8D8", x"D8D7D5D3", x"D1D2D1CC", x"C9CBCED0", x"CDC6C4C5", x"C2BEBAB4", x"AEABA7A7", x"A8A7A5A2",
									 -- x"A4A19E9C", x"9B999897", x"9B9B9895", x"94959593", x"90908F8C", x"8B8A8580", x"807F8083", x"84838385",
									 -- x"8A908F8D", x"9196989A", x"9FA3A9AD", x"AFAEADAD", x"AFB2AFB0", x"AFADB1B0", x"ADADACAB", x"ACADABA9",
									 -- x"A9A7A5A4", x"A09A9694", x"91909191", x"908F9195", x"95999A97", x"95979693", x"9B989595", x"98999895",
									 -- x"9A9F9F9E", x"A0A2A2A4", x"A29FA0A3", x"A49F9D9D", x"9E9B9898", x"98969494", x"99949399", x"9A929096",
									 -- x"97989792", x"8E8D8C8B", x"88878C88", x"85827B7C", x"77777572", x"7172716F", x"6E717271", x"71716F6C",
									 -- x"68676768", x"68666566", x"63615F5F", x"605F5E5C", x"5B565250", x"51514E4B", x"4B4B4946", x"45454341",
									 -- x"3F3D3A39", x"3A3B3936", x"36343334", x"34322F2F", x"31333332", x"31323332", x"34363838", x"36353637",
									 -- x"CCCDCECF", x"CECECECF", x"CDCDCDCE", x"CFD0D0D0", x"D0CFD0D1", x"D1D1D1D2", x"D6D6D7D8", x"D9D9D8D8",
									 -- x"D8D9D7D4", x"D5D8D8D5", x"D5D6D7D8", x"D7D6D5D3", x"D1D2D1CF", x"CAC5C1C0", x"BCB9B6B1", x"AEACAAAA",
									 -- x"A7A3A3A2", x"9E9D9B97", x"9592908F", x"8D8B8B8C", x"8A888788", x"87828181", x"7D7A7777", x"77747272",
									 -- x"72737371", x"6F6F6F6D", x"6D6D6C6C", x"6B696765", x"63615F5E", x"5E5D5C5B", x"5A5B5C5C", x"5C5B5B5B",
									 -- x"57585958", x"57565556", x"50525353", x"52515152", x"52535556", x"56555658", x"5A5B5D5E", x"5E5E5E5F",
									 -- x"5C616566", x"67686764", x"68666769", x"6B6C6F71", x"7170736F", x"71787677", x"7B7A7A7B", x"7E818282",
									 -- x"85858585", x"87888A8B", x"8D8D8D8E", x"90939595", x"97979799", x"9B9B9997", x"9A9A9896", x"9492908F",
									 -- x"908E8D8E", x"8E8D8E8F", x"8E8E9194", x"94919091", x"95929395", x"96959699", x"95969697", x"97979797",
									 -- x"97989B9F", x"A1A2A3A5", x"A5A6A7A8", x"AAACB0B2", x"B5B2B0B1", x"B2B0AEAD", x"ADACABAC", x"ACACADAE",
									 -- x"B1B3B6B9", x"BDC0C3C5", x"CDCFD2D4", x"D5D6DBE0", x"DFE2E4E4", x"E6E9EAE9", x"EBE9E7E6", x"E8EBEEF0",
									 -- x"F0F0F1F2", x"F5F7F8F8", x"F8F9FBFD", x"FEFEFDFD", x"FCFCFCFD", x"FEFEFEFD", x"FFFDFBFB", x"FCFDFDFD",
									 -- x"FBFAF8F7", x"F8F8F7F6", x"F6F6F4F2", x"F0F0EFED", x"EDECEBEB", x"EAE8E4E2", x"DEDBD8D6", x"D5D6D5D5",
									 -- x"D4D7D7D5", x"D5D6D4D1", x"D2D1CECB", x"CBCED0D0", x"CAC0BCBD", x"BCBBB7AF", x"ABA7A3A2", x"A2A19D99",
									 -- x"9C999695", x"95959390", x"96989792", x"90939390", x"8E8C8A88", x"88888480", x"7D7D7E81", x"82818182",
									 -- x"8C8F8D8A", x"8E919192", x"9A9EA4A7", x"A8A8A9AA", x"ACAEAAAB", x"ABA8ADAC", x"A6A8A8A6", x"A6A6A5A3",
									 -- x"A3A2A1A0", x"9B959292", x"928F8D8E", x"8F8E8E8F", x"93959592", x"9192918F", x"94929294", x"98999693",
									 -- x"97979A9B", x"9B9FA3A3", x"A2A0A0A2", x"A19F9FA2", x"A19D9A99", x"98969393", x"999A9699", x"9F96919D",
									 -- x"989B9D9A", x"95939292", x"8E8B8C87", x"82817B7D", x"73777978", x"76777879", x"75797B78", x"77787671",
									 -- x"6E6D6D6C", x"6A68696B", x"66666463", x"62615F5E", x"5C585353", x"5556524E", x"4D4D4C4A", x"49484644",
									 -- x"42413D3B", x"3C3E3D3A", x"39373638", x"39373635", x"36383734", x"33353535", x"393A3B3A", x"38373738",
									 -- x"CACBCCCD", x"CDCDCDCD", x"CACAC9CA", x"CBCBCAC8", x"CECBCCCF", x"CFCDCDCF", x"D2D3D4D5", x"D6D6D6D7",
									 -- x"D7D9D7D3", x"D4D9D8D3", x"D3D4D6D7", x"D7D5D4D2", x"D1D2D2CF", x"CAC6C4C3", x"C0C0BCB4", x"AEADABA8",
									 -- x"A7A3A2A2", x"9E9D9B97", x"9794918F", x"8C8A8A8B", x"88868689", x"88848386", x"817C7877", x"78777574",
									 -- x"74767673", x"706F6E6E", x"6D6C6C6D", x"6D6B6866", x"65636263", x"62605E5E", x"5E5E5E5E", x"5D5C5D5D",
									 -- x"58595958", x"57565555", x"51525354", x"53515150", x"52505155", x"5554565B", x"59595B5C", x"5D5D5C5B",
									 -- x"5C5F6160", x"60636565", x"66656667", x"68686A6D", x"6A696D6B", x"6E757577", x"79777575", x"787C7F81",
									 -- x"81818282", x"83848687", x"85888B8C", x"8E919190", x"93939394", x"96969594", x"97969695", x"93929190",
									 -- x"908D8C8C", x"8C8C8E90", x"8F919497", x"98979798", x"9C9A999A", x"9A9A9A9D", x"9A9B9C9C", x"9D9D9D9D",
									 -- x"9FA1A4A6", x"A7A7A9AB", x"ABABACAD", x"AEB1B5B7", x"BCBAB7B6", x"B6B6B4B2", x"B2B1B1B2", x"B1B0B0B2",
									 -- x"B4B7BBBE", x"C2C5C8CA", x"D5D7D9D9", x"D9DADDE0", x"E1E2E3E4", x"E6EAEBEA", x"ECEBEAEA", x"EBECEDED",
									 -- x"EFF0F0F2", x"F4F5F5F5", x"F8F9FBFC", x"FDFDFDFD", x"FCFCFCFD", x"FEFEFEFD", x"FEFDFAFA", x"FBFDFDFD",
									 -- x"FAF9F8F8", x"F8F8F7F6", x"F5F3F1F0", x"F1F2F0EE", x"ECEBEAEA", x"E9E6E2DF", x"DCD9D6D4", x"D5D6D5D5",
									 -- x"D2D6D6D2", x"D1D4D3CE", x"CFCCC9C9", x"CCCFCFCD", x"C8BFBAB9", x"B8B8B5AE", x"ABA6A09D", x"9D9D9A98",
									 -- x"96959392", x"93949391", x"92969590", x"8F92918C", x"8D8A8784", x"8483817F", x"7E7D7B7B", x"7C7E8082",
									 -- x"868A8987", x"8A8D8E90", x"979B9FA1", x"A3A6A8A9", x"ABACA7A7", x"A5A3A6A5", x"A2A4A5A3", x"A1A1A09F",
									 -- x"9E9C9B9A", x"97929090", x"928F8C8C", x"8D8C8C8D", x"8F91918F", x"8E8F8E8D", x"8A8E9294", x"93939596",
									 -- x"97959A9C", x"999DA2A0", x"A29F9EA0", x"A09E9FA0", x"9E9E9D9B", x"95919194", x"959C9B98", x"9B9C9A9C",
									 -- x"999B9B9A", x"97959493", x"908C8A83", x"7E7E797B", x"767B7F7F", x"7E7E7F81", x"7F83837E", x"7C7E7C77",
									 -- x"75757572", x"6E6B6B6C", x"6B6B6A67", x"6463615E", x"5E5B5858", x"59585552", x"51504F4D", x"4C4B4948",
									 -- x"4644413E", x"3E40403F", x"3C3B3B3C", x"3E3E3C3B", x"3D3D3C38", x"37373838", x"3B3B3B3A", x"39383838",
									 -- x"C8C9C9CA", x"CACACAC9", x"C8C8C7C8", x"C9C9C7C6", x"CBC8C8CB", x"CCC9C9CC", x"CFD0D2D3", x"D3D3D3D4",
									 -- x"D3D5D3D0", x"D1D6D4CF", x"D0D1D3D5", x"D5D5D3D2", x"D2D2D1CE", x"CBC8C7C7", x"C3C4C0B7", x"B1B0AEAA",
									 -- x"A8A4A3A2", x"9E9D9B96", x"99969391", x"8F8D8C8E", x"8B89888A", x"8A878789", x"857F7A79", x"7A797777",
									 -- x"75777672", x"6E6D6E6E", x"6B6B6B6D", x"6E6D6A67", x"66646365", x"65626060", x"61615F5D", x"5C5B5C5D",
									 -- x"5B5A5858", x"58575553", x"53535354", x"54535150", x"52505052", x"5353575C", x"57585A5C", x"5C5C5B5A",
									 -- x"5D5F5F5E", x"5E606364", x"63626264", x"63636567", x"68676B6A", x"6B706F72", x"74737373", x"75787B7C",
									 -- x"7C7D7F7F", x"80808283", x"82868A8A", x"8A8B8D8E", x"8E8F9192", x"92929293", x"92929191", x"90908F8F",
									 -- x"918F8D8D", x"8E8E9092", x"9596989C", x"9D9D9D9F", x"A1A09F9F", x"9F9E9FA0", x"A0A0A1A2", x"A2A3A3A3",
									 -- x"A5A7A9A9", x"AAACAEB0", x"AFAFB0B1", x"B3B7BBBE", x"C3C0BDBB", x"BBBBBAB8", x"B6B5B5B6", x"B5B4B3B4",
									 -- x"B7BCC1C5", x"C7CACFD3", x"DADCDDDD", x"DCDDDFE1", x"E2E2E3E3", x"E6E9E9E9", x"E9EAEBEC", x"EDEDEBE9",
									 -- x"EDEEEFF0", x"F2F4F4F4", x"F8F9FAFB", x"FBFCFDFE", x"FCFCFCFD", x"FEFEFEFD", x"FDFBFAFA", x"FBFCFCFB",
									 -- x"F9F9F8F8", x"F8F8F6F6", x"F4F1EFEF", x"F0F1F0EE", x"EBEAE9E8", x"E7E4E0DC", x"DAD7D4D4", x"D5D6D5D4",
									 -- x"D2D6D5D1", x"D0D2D1CC", x"CDCAC8CA", x"CCCDCBC9", x"CBC4C0BC", x"B7B6B4AF", x"AAA59F9B", x"9A999795",
									 -- x"96969592", x"90929291", x"8F92928F", x"8E8F8B85", x"89868584", x"84817E7B", x"7D7C7977", x"787B7E80",
									 -- x"7C828485", x"898C8F94", x"95989A9C", x"A1A6A9A8", x"A8A9A2A2", x"A09EA1A0", x"A0A2A29F", x"9E9D9C9B",
									 -- x"9B979494", x"93908E8D", x"8D8B8A8A", x"8B8C8E91", x"8B8D8E8E", x"8D8D8C8B", x"878B8F90", x"8F909294",
									 -- x"9593999D", x"999A9E9C", x"9E9C9B9D", x"A0A09F9F", x"9C9C9C9A", x"95929396", x"92949A9C", x"9A9FA5A0",
									 -- x"A09D9A99", x"97949190", x"908B8A83", x"80817D7F", x"85878B8D", x"8C8B8B8B", x"8D8F8C84", x"8182817C",
									 -- x"7A7C7B77", x"726F6E6E", x"70706E6A", x"67666461", x"605F5F5D", x"5B595857", x"55535150", x"4E4D4C4C",
									 -- x"48474441", x"41434342", x"3F3F3E3E", x"3F3F3D3B", x"3E3F3E3B", x"3A3A3B3B", x"3C3C3B3A", x"39383939",
									 -- x"CAC9C9C9", x"CAC9C8C7", x"C6C6C6C6", x"C7C7C7C6", x"C6C5C4C5", x"C5C5C6C7", x"CBCCCECF", x"CFCFCFD0",
									 -- x"D0D1D1CF", x"D0D2D1CD", x"CCCDCFD1", x"D2D2D2D1", x"D2D1CFCC", x"CBC9C8C8", x"C2C2BFBA", x"B6B4B2AE",
									 -- x"AAA6A5A4", x"A09E9C97", x"99969493", x"918E8E8F", x"8D8B8A89", x"8A898887", x"86817C7B", x"7B7A7979",
									 -- x"77787671", x"6D6C6D6D", x"6B6B6B6C", x"6C6C6A69", x"65636366", x"66636162", x"61605F5C", x"5A595A5A",
									 -- x"5D5B5858", x"59595754", x"55545454", x"54545250", x"52515050", x"50515559", x"5557595B", x"5B5B5B5B",
									 -- x"5E5F5F5F", x"5E5E5F5F", x"62606061", x"61616263", x"65646967", x"686C6A6D", x"6C6E7174", x"76777777",
									 -- x"7A7C7E7E", x"7E7E8081", x"83858687", x"8585898F", x"898C8E90", x"90909294", x"92929191", x"90909090",
									 -- x"95929191", x"92939598", x"9A9A9C9F", x"9F9FA0A2", x"A5A4A4A4", x"A4A5A5A6", x"A6A7A8A8", x"A9AAAAAA",
									 -- x"A9ABACAC", x"ADB0B3B4", x"B3B4B5B6", x"B9BDC1C4", x"C7C5C1BE", x"BFC1C0BF", x"BBBABABB", x"BBB9B9BA",
									 -- x"BBC0C6C9", x"CACDD3D8", x"DBDEE0E0", x"E0E1E3E3", x"E3E2E2E3", x"E5E7E7E6", x"E6E7E9EB", x"ECEBE9E7",
									 -- x"EAEAECEE", x"F1F3F4F4", x"F6F8F9FA", x"FAFBFDFE", x"FCFCFCFC", x"FDFEFEFD", x"FCFBFAFB", x"FCFCFAF9",
									 -- x"F9F9F9F8", x"F8F7F6F6", x"F4F0EDED", x"EEEDECEC", x"EBEAE8E7", x"E6E3DEDB", x"D9D6D4D4", x"D6D7D5D3",
									 -- x"D2D5D4D1", x"D0D0CFCB", x"CDCBCACB", x"CCCBC8C7", x"CEC9C5BF", x"B7B4B3AE", x"A8A5A19D", x"99969492",
									 -- x"989A9993", x"9090908E", x"8E8E8D8D", x"8D8B857F", x"83828284", x"84817B78", x"79797876", x"7678797A",
									 -- x"787F8283", x"86878A90", x"9195989A", x"9FA5A7A5", x"A2A29C9D", x"9D9B9F9C", x"9E9E9D9A", x"99999896",
									 -- x"96928E8E", x"8F8D8B8A", x"8B8A8A8A", x"89898B8E", x"88898B8B", x"8A8A8989", x"8988888A", x"8D8E8E8D",
									 -- x"8E8F959B", x"9B9C9E9E", x"9D9B9A9C", x"9F9F9D9A", x"9C989697", x"98979696", x"968E97A1", x"9D9EA4A3",
									 -- x"A19C9795", x"9593908F", x"8C888985", x"85888587", x"8B8D9195", x"98989798", x"9A979189", x"8382817F",
									 -- x"7B7C7C79", x"76747271", x"7374716D", x"6B6B6966", x"64656562", x"5F5C5C5C", x"58565352", x"51504F50",
									 -- x"4A494744", x"44464645", x"4242413F", x"3F3F3D3A", x"3D3F3F3E", x"3D3E3E3E", x"3E3D3C3B", x"3A3A3B3B",
									 -- x"C9C9C8C9", x"C9C9C7C6", x"C4C4C4C3", x"C2C2C2C3", x"C3C3C1BF", x"BFC1C3C4", x"C5C7C9CA", x"C9C9CBCC",
									 -- x"CDCECECE", x"CECECDCC", x"CACBCDCE", x"CECECECD", x"CFCDCAC9", x"C9C8C6C4", x"C1C0BDBB", x"B9B7B4B1",
									 -- x"ACA8A7A6", x"A2A09F9A", x"9A979594", x"928F8E8F", x"8C8D8B89", x"8B8E8B85", x"85817E7D", x"7C797979",
									 -- x"78787670", x"6C6B6A6A", x"6A6A6A6A", x"69686869", x"67646467", x"67636263", x"6161615F", x"5D5B5B5A",
									 -- x"5D5B5A5A", x"5A5A5958", x"57575756", x"55535352", x"52535250", x"4F515456", x"5456595A", x"59595A5B",
									 -- x"5E5E5D5D", x"5E5D5D5C", x"615F5E60", x"61616162", x"62616564", x"6568676B", x"686A6E71", x"74757677",
									 -- x"78797A7A", x"7A7A7D7F", x"827F8084", x"8483878E", x"88898C8E", x"8F909192", x"95949392", x"92939495",
									 -- x"97959495", x"97989B9E", x"9F9FA1A3", x"A4A3A4A6", x"A9A9AAAA", x"AAABACAC", x"ACADAFB1", x"B2B2B1B1",
									 -- x"B0B1B1B1", x"B3B7B8B7", x"B9B9BABB", x"BDC0C3C6", x"C7C5C2BF", x"C0C3C4C2", x"C1BFC0C1", x"C2C1C2C4",
									 -- x"C3C6CACD", x"CFD2D7DB", x"DEE2E4E4", x"E4E6E6E5", x"E4E3E2E3", x"E4E5E4E3", x"E5E4E5E6", x"E7E7E7E6",
									 -- x"E8E8E9EB", x"EEF0F2F2", x"F4F6F9FA", x"FAFAFCFE", x"FCFCFBFC", x"FDFEFEFD", x"FDFCFBFB", x"FBFBFAF9",
									 -- x"F9F9F8F7", x"F6F5F4F4", x"F3EFECEC", x"EBEAE9E9", x"E9E8E6E5", x"E3E1DDDA", x"D8D6D4D5", x"D7D7D4D1",
									 -- x"D2D2D2D0", x"CFCDCBCA", x"C9C9C9CB", x"CBC9C8C9", x"CECAC6C0", x"B8B5B3AD", x"A9A8A5A0", x"9B989798",
									 -- x"9A9C9B97", x"9596948F", x"8E8A878A", x"8D8A8480", x"807D7C7E", x"7F7C7977", x"75767572", x"72747474",
									 -- x"767B7D7E", x"81818185", x"8B91989B", x"9EA2A29F", x"9C9D9799", x"99989C9A", x"9A999794", x"93949290",
									 -- x"908D8A8A", x"89888889", x"88878889", x"88868687", x"85868686", x"85858585", x"86858586", x"898A8B8A",
									 -- x"898D9196", x"9A99999D", x"9A9A999A", x"9B9B9997", x"9A979596", x"97979696", x"9894989F", x"9F9D9D9D",
									 -- x"9C989392", x"918F8E8E", x"89868A89", x"8B908D8F", x"8C8F949B", x"9E9F9FA1", x"9F9A928C", x"87828283",
									 -- x"7E7F7E7B", x"7A7B7B79", x"7978746F", x"6E706D69", x"69696866", x"63616060", x"5A575555", x"55525152",
									 -- x"4B4B4A48", x"47484846", x"45454442", x"4243413E", x"40424342", x"42424140", x"42403E3D", x"3D3D3E3E",
									 -- x"C5C5C5C5", x"C7C7C6C4", x"C2C3C2C0", x"BDBCBDBE", x"C1C2C0BC", x"BCC0C3C2", x"C0C2C5C6", x"C6C6C7C9",
									 -- x"CAC9CBCC", x"CBC9C8C9", x"CBCBCCCC", x"CBCAC9C9", x"CBC8C6C7", x"C8C7C4C0", x"C1BEBCBC", x"BBB8B3B1",
									 -- x"ADA9A9A8", x"A4A2A19C", x"9E9B9997", x"94908E8E", x"8C8E8D8C", x"90959188", x"83817F7E", x"7C797879",
									 -- x"78787570", x"6B6A6866", x"68696967", x"65646567", x"69656568", x"68646365", x"63646464", x"625F5D5D",
									 -- x"5B5C5C5B", x"5A5A5B5B", x"595B5B59", x"55535355", x"50545451", x"50545555", x"55585A5A", x"58575859",
									 -- x"5E5C5A5A", x"5C5C5D5D", x"5F5C5B5E", x"60616060", x"64626563", x"62656368", x"68696B6D", x"70737779",
									 -- x"73747574", x"7374787A", x"7D797B84", x"8784858C", x"89898A8D", x"8F91908E", x"94949392", x"93949697",
									 -- x"97959597", x"999B9EA1", x"A3A3A6A9", x"ABAAABAD", x"ADAEAFAE", x"AFAFAFAF", x"B0B2B5B7", x"B8B7B6B5",
									 -- x"B7B8B7B7", x"B9BCBCB9", x"BEBEBEBE", x"BEBFC2C3", x"C6C4C0BE", x"BFC3C5C3", x"C5C4C4C6", x"C7C8C9CB",
									 -- x"CDCECFD2", x"D4D8DBDD", x"E1E5E8E8", x"E7E8E8E5", x"E5E3E2E3", x"E4E4E2E1", x"E5E3E2E1", x"E2E4E6E6",
									 -- x"E7E7E8EA", x"ECEEEFEF", x"F2F5F8FA", x"FAFAFCFD", x"FDFCFBFB", x"FCFDFEFE", x"FFFDFBFB", x"FBFBFAF9",
									 -- x"F7F7F6F5", x"F3F2F2F2", x"F1EEEBEB", x"EAE8E7E9", x"E7E5E3E2", x"E1DFDCD9", x"D8D6D4D5", x"D8D7D4D1",
									 -- x"D0CFCECF", x"CDCAC7C7", x"C5C5C7CA", x"C9C8CACD", x"CECAC7C1", x"BBB9B7B0", x"ADABA7A1", x"9C9B9EA1",
									 -- x"999B9C9B", x"9C9E9B94", x"8E868389", x"8E8C8784", x"827C7776", x"76757677", x"7474726E", x"6D707271",
									 -- x"6F737578", x"7E7F7E80", x"858F989B", x"9D9F9D9A", x"999A9596", x"97969997", x"9795928F", x"8F908E8B",
									 -- x"8B898887", x"85848588", x"82828488", x"89878584", x"84838382", x"81808182", x"7E828686", x"8585898C",
									 -- x"898E8F91", x"95918D93", x"93949697", x"98999999", x"97989897", x"93909295", x"929C9A96", x"9EA09998",
									 -- x"9D999592", x"8E8A898B", x"8A888D8E", x"92969395", x"95979DA2", x"A3A2A3A6", x"A29B9491", x"8C86868A",
									 -- x"84848280", x"80838382", x"7D7C7771", x"70726F6A", x"6C6B6968", x"66656463", x"5B585758", x"57545253",
									 -- x"4B4D4C4A", x"4A4A4947", x"47484746", x"48494845", x"44474847", x"46454341", x"45444140", x"3F404041",
									 -- x"C7C5C3C3", x"C4C4C2C1", x"C0BFBDBC", x"BCBCBCBC", x"BDBDBDBC", x"BCBCBDBD", x"BDBEC0C3", x"C4C3C2C1",
									 -- x"C4C6C8C8", x"C8C7C7C7", x"C7C9C8C6", x"C7C5C4C6", x"C4C5C6C4", x"C0BEBFC1", x"BDBEBCB9", x"B6B5B3B0",
									 -- x"AEACAAA7", x"A3A1A1A1", x"9B9A999A", x"97928F8F", x"918E8D8F", x"8F8D8B8B", x"81828280", x"7E7D7A76",
									 -- x"7B78736F", x"6D6C6966", x"69686765", x"64646565", x"63646566", x"66656363", x"64636160", x"60616262",
									 -- x"595A5C5D", x"5C5A5A5C", x"5D5B5856", x"56575959", x"59565454", x"54545659", x"555A5C58", x"55585B5C",
									 -- x"59595958", x"57585A5B", x"5C5B5B5D", x"6061605F", x"62616060", x"63666561", x"656B6C6A", x"6B71726F",
									 -- x"73717071", x"72737475", x"797D8182", x"82838689", x"88898789", x"8F918F90", x"94959596", x"96969595",
									 -- x"9396999A", x"9C9FA3A6", x"A9AAABAD", x"AFB1B3B5", x"B5B4B3B3", x"B4B6B8BA", x"BEBDBCBD", x"BEBFBEBD",
									 -- x"BDC1BFBC", x"BDBEBEC1", x"C3C1BFC1", x"C3C4C3C1", x"C5C4C4C4", x"C5C7C8C9", x"C9CACBCA", x"CACBCED0",
									 -- x"D1D2D4D7", x"DADCDEDF", x"E3E5E6E7", x"E8EAE8E5", x"E6E3E1E2", x"E4E5E3E1", x"E1E1E1E1", x"E2E3E5E6",
									 -- x"E6E5E7EA", x"ECECEEF1", x"F1F6F6F7", x"F9F9F9FD", x"FDFCFCFD", x"FDFEFEFF", x"FCFBFAFA", x"FBFBFAF9",
									 -- x"F5F5F5F5", x"F4F4F2F1", x"EEEBE8E7", x"E8E9E8E6", x"E5E3E1E0", x"DEDBD9D7", x"D8D5D3D5", x"D6D4D1CF",
									 -- x"D0CCCCCD", x"C8C7C9C9", x"C3C5C7C7", x"CACECFCD", x"CECECDC6", x"BEB6B3B3", x"ACAEAA9F", x"9DA5AAA8",
									 -- x"A4A19FA0", x"9E9A9899", x"93868084", x"84838383", x"7C787675", x"73717377", x"6C6E6D6A", x"696C6E6D",
									 -- x"6B717374", x"77777B82", x"828A9399", x"9B9B9894", x"95918D8D", x"91949594", x"93909190", x"8C8C8E8C",
									 -- x"88868584", x"807D7F83", x"7E808282", x"83848380", x"8382817E", x"7A7A7C7E", x"7C7F807F", x"80838483",
									 -- x"87878A90", x"9392908F", x"93929193", x"9595928F", x"96939293", x"918D8F95", x"97949397", x"98959596",
									 -- x"9597928A", x"8B908D85", x"898B8F92", x"96989999", x"97A0A8AB", x"ABACA9A4", x"A39D9793", x"908B8887",
									 -- x"85848688", x"888A8A85", x"807E7A74", x"7475726C", x"70706F6B", x"69686665", x"625D595A", x"5A575452",
									 -- x"5252504E", x"4D4F4F4D", x"49494A4A", x"4A494746", x"48484949", x"48454444", x"45444548", x"46424246",
									 -- x"C9C8C7C5", x"C3C2C0C0", x"BDBCBBBA", x"BABAB9B9", x"BBBABAB9", x"B9BABABB", x"BBBCBEC0", x"C0C0BFBF",
									 -- x"C1C2C2C3", x"C4C4C4C4", x"C3C5C4C3", x"C5C3C1C2", x"C4C3C1BE", x"BBBBBDBF", x"BCBCBCB9", x"B6B4B1AE",
									 -- x"AAA9A7A5", x"A29F9E9D", x"9B9A9999", x"97939191", x"93908F91", x"908D8B8A", x"85858481", x"807F7C7A",
									 -- x"7976726E", x"6C6A6867", x"68686665", x"65656565", x"67666666", x"66656565", x"64636160", x"60606061",
									 -- x"5E5D5D5F", x"5F5D5B5B", x"5B5B5B5C", x"5C5B5A59", x"5B585656", x"55545557", x"585A5A58", x"58595A5B",
									 -- x"59595958", x"57575859", x"5B5B5C5E", x"60605F5D", x"5F606162", x"63636464", x"64676766", x"686D7171",
									 -- x"75737375", x"76757677", x"777A7F81", x"81828587", x"8A8B8A8C", x"92949294", x"9697999A", x"9A9A9A99",
									 -- x"989B9EA1", x"A2A4A7A9", x"AAADB1B5", x"B8B9B9B9", x"BDBCBCBC", x"BDBEBFBF", x"C1C1C1C2", x"C4C4C4C4",
									 -- x"C2C5C2C0", x"C1C1C1C5", x"C6C6C7C6", x"C5C5C4C4", x"C7C7C7C7", x"C8CACDD0", x"CDCECFCF", x"D0D1D4D6",
									 -- x"D9D9DADB", x"DDE0E2E3", x"E5E6E7E8", x"E9EAE9E6", x"E7E4E2E3", x"E5E5E3E1", x"DEDEDFDF", x"E0E2E3E3",
									 -- x"E5E4E6E8", x"EAEBEEF2", x"F2F5F4F5", x"FAFBFAFD", x"FDFDFDFC", x"FCFCFCFC", x"FAFAF9F9", x"FBFBFAFA",
									 -- x"F5F5F4F3", x"F3F2F1F0", x"EFECE9E7", x"E8E8E7E5", x"E3E2E0DE", x"DCDAD8D7", x"D6D3D1D1", x"D1CECCCB",
									 -- x"D0CCCBCB", x"C6C4C5C5", x"C2C4C5C6", x"C9CCCDCC", x"CBC9C6C1", x"BCB6B1AE", x"ADADA8A2", x"A3A9ABA7",
									 -- x"9F9D9D9F", x"9F9B9897", x"90878382", x"7F7F8283", x"79777675", x"73716F70", x"6B686667", x"66646669",
									 -- x"6A6F7071", x"74767980", x"848C9397", x"9795928F", x"8C8B8B8F", x"94969390", x"908B8A8A", x"898A8A86",
									 -- x"8582807F", x"7E7C7D7F", x"7B7E7F7F", x"8081807D", x"787A7C7C", x"7B7A797A", x"7A7C7C7B", x"7B7F8181",
									 -- x"8383868B", x"8D8D8D8D", x"91919292", x"91908F8E", x"8F91928F", x"8D8E8F90", x"928E8D90", x"918F9092",
									 -- x"9495938D", x"8C8F8D88", x"8E929597", x"9A9EA0A0", x"A5AAADAF", x"B0AFA8A0", x"A6A09A97", x"948F8C8B",
									 -- x"8B88888A", x"8A8D8C86", x"82807C77", x"75757574", x"75767470", x"6D6C6A69", x"67625E5E", x"5F5C5957",
									 -- x"56555350", x"5051504E", x"4C4D4E4F", x"4F4E4E4E", x"4E4D4D4E", x"4C484748", x"47464749", x"48444448",
									 -- x"CCCCCBC8", x"C3C0BFBE", x"BCBBB9B9", x"B8B8B7B7", x"B7B6B5B5", x"B5B6B7B7", x"B7B8B9BA", x"BBBCBCBB",
									 -- x"BDBCBBBC", x"BEC0C0C0", x"C1C3C1C1", x"C4C1BDBD", x"BEBCBAB8", x"B7B8B9BA", x"B9BBBAB8", x"B5B3B0AD",
									 -- x"AAA9A8A6", x"A3A19E9D", x"9C9B9A99", x"98959393", x"918F8F90", x"908D8987", x"8484827F", x"7D7C7B7A",
									 -- x"7775726E", x"6B6A6969", x"66656565", x"65656464", x"68676564", x"64646565", x"64646362", x"61616161",
									 -- x"64616062", x"62605D5C", x"5C5C5D5E", x"5E5D5C5B", x"5C5A5858", x"57555557", x"5B59595A", x"5A59595A",
									 -- x"595A5A59", x"58575757", x"58595C5E", x"5F5F5E5D", x"5E5F6264", x"62606267", x"67676767", x"686A6D6F",
									 -- x"71717376", x"77757576", x"777A7E81", x"83858687", x"8B8E8E90", x"95969699", x"9B9C9D9F", x"9F9F9E9D",
									 -- x"9C9FA3A5", x"A6A8AAAC", x"AFB2B7BB", x"BEBFBFBE", x"C1C1C2C3", x"C3C4C3C3", x"C4C4C5C6", x"C8C9C9C9",
									 -- x"C7C7C4C3", x"C4C2C3CA", x"CBCED0CE", x"CAC7C8CA", x"CCCBCBCA", x"CBCED2D4", x"D1D3D4D6", x"D7D8DBDE",
									 -- x"DFDFDEDF", x"E0E3E5E7", x"E8E9E9E9", x"E9EBE9E7", x"E8E6E4E4", x"E5E5E3E1", x"DDDDDEDF", x"E0E0E1E1",
									 -- x"E3E3E4E6", x"E7E9EDF0", x"F2F4F3F5", x"FBFDFCFD", x"FEFDFDFC", x"FBFAFAFA", x"FAFAF9F9", x"FAFAF9F9",
									 -- x"F5F4F3F2", x"F1F1F0EF", x"EEEBE8E7", x"E7E7E6E4", x"E2E1DFDC", x"DAD8D5D4", x"D5D2D0CE", x"CDCBCBCC",
									 -- x"D1CDCDCC", x"C6C4C5C4", x"C2C3C3C4", x"C6C9CBCA", x"C9C5C1BE", x"BCB9B4AF", x"B0ABA6A5", x"AAAEAAA5",
									 -- x"9C9C9D9F", x"A09C9794", x"8B878480", x"7A7B8081", x"77777471", x"706F6C68", x"6B626065", x"645E5F67",
									 -- x"6A6D6D6E", x"7275777D", x"7E858D8F", x"8F8E8C8A", x"8B888688", x"8E91908E", x"8E888687", x"8788857E",
									 -- x"7E7A7778", x"79787878", x"78797B7B", x"7B7C7B79", x"75767879", x"78777473", x"787A7B7B", x"7C7E7F7F",
									 -- x"82828487", x"89898A8D", x"8E909190", x"8D8A8A8B", x"848B8D87", x"868C8D88", x"8C898789", x"8A898B8D",
									 -- x"8E909190", x"8F909190", x"90979B9C", x"9FA6A9A8", x"B0B4B7B6", x"B5B2ADA7", x"A5A19D9B", x"99969393",
									 -- x"95908F90", x"9195938B", x"8784807C", x"7876787B", x"797A7975", x"71706E6D", x"6B666262", x"62605D5B",
									 -- x"5B595654", x"54565350", x"53545454", x"52505051", x"51504F4F", x"4C494849", x"4948494B", x"4A464749",
									 -- x"CECECCC9", x"C5C2BFBD", x"BDBCB9B8", x"B7B6B6B5", x"B4B3B2B1", x"B1B2B3B4", x"B3B4B5B5", x"B5B7B7B7",
									 -- x"BAB8B6B7", x"BABDBEBE", x"C0C1BFBE", x"C1BEB8B6", x"B4B4B4B5", x"B6B6B5B4", x"B7B8B8B5", x"B4B3B1AE",
									 -- x"ACAAA9A7", x"A5A2A09F", x"9D9C9A99", x"97959393", x"8E8E8F90", x"908E8A87", x"8282807D", x"7A7A7977",
									 -- x"7776736E", x"6B696969", x"65666667", x"67666666", x"68676664", x"64646465", x"65656564", x"64636363",
									 -- x"66646364", x"64615F5E", x"5E5E5D5B", x"5B5B5C5D", x"5C5B5A59", x"59585858", x"5B58595B", x"5C59595B",
									 -- x"5A5A5B5B", x"5A595858", x"56585A5C", x"5D5E5F5F", x"605F6264", x"625E6169", x"68686A6D", x"6D6C6C6E",
									 -- x"6F6E7074", x"76747577", x"7B7C7E82", x"86898B8C", x"8C919293", x"9798999D", x"9EA0A1A2", x"A2A1A09F",
									 -- x"9FA2A6A8", x"A9ABAEB1", x"B7B8BABC", x"BEC0C2C3", x"C3C3C4C5", x"C6C7C7C7", x"C7C8CACC", x"CDCECECE",
									 -- x"CCC9C6C6", x"C7C4C6CF", x"D2D5D7D4", x"CECBCDD0", x"D1CFCDCD", x"CFD2D3D4", x"D5D7D9DA", x"DBDDE0E3",
									 -- x"E1E1E2E3", x"E5E7E9EB", x"EAEBEBE9", x"E9EAEAE8", x"E9E8E6E6", x"E6E5E4E3", x"DFDFDFDF", x"DFE0E1E2",
									 -- x"E2E2E3E5", x"E6E8EBED", x"F1F4F4F7", x"FCFDFCFE", x"FEFEFDFC", x"FBFAF9F9", x"FBFAFAF9", x"F8F7F6F6",
									 -- x"F5F4F2F0", x"F0EFEFEE", x"EAE8E6E5", x"E5E5E5E3", x"E3E1DEDB", x"D8D5D2D0", x"D2D0CECC", x"CBCACCD0",
									 -- x"CECBCCCB", x"C6C5C6C4", x"C3C3C3C3", x"C5C6C7C6", x"C7C2BDBB", x"BBBAB6B3", x"B2ABA5A7", x"ADADA8A3",
									 -- x"9E9D9D9F", x"9F9B9590", x"8785827D", x"797C7F7C", x"7675716B", x"6A6B6964", x"675F5C61", x"605B5C63",
									 -- x"686C6C6C", x"71747579", x"777E8689", x"89888786", x"87838081", x"878B8C8B", x"8E888686", x"8584817A",
									 -- x"78767373", x"74747474", x"73757777", x"77777777", x"76757474", x"74747473", x"76787B7D", x"7E7D7C7C",
									 -- x"82828385", x"85848689", x"888A8C8B", x"87848383", x"83898A86", x"868C8D89", x"89878687", x"8887898B",
									 -- x"8C8D8F91", x"91919295", x"939BA0A1", x"A5AEB4B3", x"B7BFC4C0", x"B8B3B1B1", x"AAA7A4A1", x"9F9C9A99",
									 -- x"99969697", x"97999790", x"8C878381", x"7E7A7B7F", x"7A7C7B77", x"74727270", x"6F6B6765", x"64625F5D",
									 -- x"5E5C5857", x"595B5854", x"58595957", x"55535354", x"53514F4E", x"4B494A4C", x"4C4B4C4D", x"4B49484A",
									 -- x"CFCDCBCA", x"C8C5C0BD", x"BEBCB8B6", x"B4B4B4B4", x"B1B0AFAE", x"ADAEAFB0", x"AEB0B0AF", x"B0B2B3B2",
									 -- x"B7B5B3B4", x"B7BABCBC", x"BBBCBABA", x"BCB8B2B0", x"B0AFB0B1", x"B3B3B1AF", x"B4B5B5B3", x"B2B2B2B0",
									 -- x"ACAAA7A4", x"A3A2A09F", x"9E9D9B97", x"95939290", x"8F909091", x"918F8A87", x"8384827E", x"7B7A7977",
									 -- x"7775726D", x"6A686868", x"67686969", x"6A696968", x"69696867", x"67666666", x"65656566", x"66666565",
									 -- x"65656566", x"64616061", x"605F5D5A", x"59595B5D", x"5C5C5B5A", x"5A5A5959", x"5A585A5D", x"5C595A5E",
									 -- x"5A5A5B5C", x"5D5D5C5B", x"5A5A5B5C", x"5C5E6061", x"63606063", x"6361646C", x"66676A6E", x"70707274",
									 -- x"73727377", x"7875777B", x"7D7D7F83", x"888C8F90", x"8E939495", x"999A9BA0", x"A0A1A3A4", x"A4A3A2A1",
									 -- x"A5A7A9AA", x"ACAFB4B8", x"BDBDBEBF", x"C2C4C7C8", x"CACACACA", x"CBCCCDCD", x"CDCFD1D3", x"D4D4D3D3",
									 -- x"D1CECACB", x"CCC9CBD5", x"D8D9D9D6", x"D3D1D3D5", x"D6D2CFD0", x"D4D7D6D4", x"D7D9DCDD", x"DEE0E3E5",
									 -- x"E5E6E7E8", x"E9EBECED", x"EBECEBE9", x"E8E9EAE9", x"EBEAE8E7", x"E6E5E5E5", x"E2E1E0DF", x"E0E1E2E3",
									 -- x"E2E4E6E7", x"E8E9EAEB", x"EFF5F7F9", x"FDFDFBFE", x"FEFDFDFC", x"FBFAFAF9", x"FAFAF9F8", x"F6F5F4F4",
									 -- x"F4F3F1EF", x"EFEEEDED", x"E9E8E6E5", x"E5E4E3E2", x"E1DFDCD8", x"D5D2D0CE", x"CDCBC9C8", x"C6C6CACE",
									 -- x"C8C6C7C7", x"C4C4C6C4", x"C4C3C2C2", x"C3C2C1C1", x"C2BEB9B5", x"B4B4B2B1", x"B2ABA6A7", x"AAA8A4A1",
									 -- x"9C9C9C9B", x"9B97928D", x"86827F7C", x"7B7F7E76", x"73726D67", x"66676560", x"605C5A5A", x"5A595A5C",
									 -- x"63696969", x"6E727376", x"767D8486", x"85848280", x"7C7B7C80", x"86888785", x"8A868585", x"817F7C77",
									 -- x"75747372", x"72727373", x"70727375", x"75747576", x"73717071", x"72747676", x"74747679", x"7A78787A",
									 -- x"7D7E8082", x"81808285", x"83848585", x"84817D7B", x"80818282", x"83858788", x"86868789", x"8989898A",
									 -- x"8F8E8E91", x"91919294", x"9BA1A6A7", x"ADB7BDBE", x"C3C9CCC7", x"BEB7B6B7", x"B5B3AFAA", x"A6A3A09E",
									 -- x"9C9B9C9C", x"98989691", x"8F8A8686", x"85818082", x"7C7D7C79", x"77777674", x"75726E6B", x"6866625F",
									 -- x"5F5D5B5A", x"5D5F5D59", x"595A5B5B", x"5A595A5B", x"57555250", x"4E4D4F51", x"4F4E4E4E", x"4D4B4A4A",
									 -- x"CFCDCBCA", x"C9C7C1BD", x"BCBAB6B3", x"B1B1B1B1", x"AEADACAB", x"AAAAABAB", x"A9ACACAA", x"ABAEAEAC",
									 -- x"B2B1B0B1", x"B3B6B8B8", x"B6B9B8B8", x"BAB6B0AF", x"B0AFAEAE", x"AEAFAEAD", x"B0B2B2B1", x"B1B2B1B0",
									 -- x"ADAAA7A4", x"A4A3A1A0", x"9E9E9B98", x"95949291", x"91919190", x"8F8D8985", x"84858480", x"7B7A7877",
									 -- x"7674706B", x"68676767", x"67676868", x"69686868", x"68686868", x"67676665", x"64646566", x"66666666",
									 -- x"64646666", x"63606062", x"5E5F5F5D", x"5B5A5B5C", x"5D5D5D5B", x"5A5B5B59", x"5A5B5C5D", x"5C5B5D5F",
									 -- x"5B5C5D5F", x"61626161", x"6362605E", x"5E5F6162", x"64626264", x"66676A6F", x"696A6C6D", x"6F727577",
									 -- x"7A78787B", x"7B77797E", x"7E7E8084", x"898D9092", x"92979899", x"9D9E9FA3", x"A1A2A4A6", x"A7A7A7A7",
									 -- x"A9AAABAC", x"ADB1B8BC", x"BFC1C3C7", x"CACDCECF", x"D3D2D1D0", x"D0D0D1D2", x"D1D3D6D8", x"D8D7D7D6",
									 -- x"D4D2CECD", x"CECCCFD7", x"DBDBDBD9", x"D7D6D8D9", x"D9D5D2D3", x"D8DBDAD8", x"DADCDFE0", x"E1E3E5E7",
									 -- x"E9E9EAEA", x"EBEBEBEB", x"ECEDECE9", x"E8E9EAEA", x"ECEBEAE8", x"E6E5E6E7", x"E4E4E2E1", x"E1E1E2E2",
									 -- x"E4E7E9E9", x"EAEBEBEB", x"EEF4F7F9", x"FCFCFBFE", x"FEFDFCFB", x"FAFAF9F9", x"F7F8F7F6", x"F5F4F3F4",
									 -- x"F1F0EFEE", x"EEEDECEB", x"EBEAE8E6", x"E4E3E1E0", x"DDDBD8D5", x"D3D1CFCE", x"CBC9C7C5", x"C3C3C6C9",
									 -- x"C3C3C5C5", x"C2C3C5C3", x"C3C1C0C1", x"C0BDBBBB", x"BEBBB6B2", x"AFADACAB", x"AEA9A5A4", x"A4A29F9D",
									 -- x"96979795", x"93918E8A", x"86807C7B", x"7C7F7B72", x"6F6E6B67", x"6563605C", x"5C5C5A57", x"585B5C59",
									 -- x"5F656665", x"6A6E7073", x"71777C7F", x"7F7F7E7C", x"7C7C7C7E", x"80828281", x"82808180", x"7B797875",
									 -- x"7071716F", x"6F707070", x"6F707274", x"73727375", x"6F707070", x"71727273", x"75727275", x"7574767B",
									 -- x"7B7B7D7F", x"807F8082", x"81818182", x"84827E79", x"7D7A7A7E", x"807E8084", x"8284888B", x"8D8D8E8F",
									 -- x"91909192", x"9495989B", x"A2A5A8AC", x"B4BDC3C5", x"CDCCCBC9", x"C7C5C1BE", x"BBBAB6B1", x"AEACAAA8",
									 -- x"A6A5A6A2", x"9C999792", x"908E8C8C", x"8C898786", x"81807F7D", x"7E7F7D7A", x"7977736F", x"6B696561",
									 -- x"61605F5F", x"6164625F", x"5E5E5E5E", x"5D5C5B5B", x"59575655", x"53525355", x"52525151", x"504E4D4C",
									 -- x"CFCECDCC", x"C9C5C1BD", x"B9B7B4B2", x"B1B0AFAF", x"ABAAA9A7", x"A6A6A6A6", x"A5A8A8A6", x"A7AAAAA7",
									 -- x"ABACACAD", x"AFB0B2B3", x"B5B8B8B7", x"B8B5B0AF", x"AEAEADAD", x"ACACABAA", x"ACAEB0B0", x"B0B0AFAC",
									 -- x"AEACA9A7", x"A7A6A4A2", x"A0A09F9C", x"9A9A9896", x"93939290", x"8F8E8B87", x"8687857F", x"7A787878",
									 -- x"77736F6B", x"69696867", x"66666767", x"67676767", x"67676767", x"67666665", x"65656767", x"68676666",
									 -- x"65646465", x"64616060", x"5D5E5F5E", x"5C5A5A5B", x"5C5D5C5A", x"5A5C5D5B", x"5D5E5E5D", x"5D5F605F",
									 -- x"60606264", x"67686868", x"6C696663", x"63646565", x"65666869", x"696B6F71", x"6F727372", x"73777A79",
									 -- x"7E7C7D80", x"7F7B7D83", x"8183868A", x"8D909293", x"989C9C9E", x"A2A3A4A7", x"A5A6A8AA", x"ACACADAD",
									 -- x"ADAEAEAE", x"B0B4BABF", x"C0C3C6CB", x"CFD2D4D5", x"D8D7D5D4", x"D3D3D4D4", x"D3D6DADB", x"DCDBDADA",
									 -- x"D6D6D2CE", x"CECFD0D6", x"DBDDDEDD", x"DBDADBDC", x"DDD9D6D5", x"D8DBDCDC", x"DEE0E2E4", x"E6E7E9EB",
									 -- x"EDECEBEB", x"EAEAEAEA", x"EDEEECE9", x"E7E9EBEC", x"EDECEBE8", x"E5E5E8EA", x"E7E7E7E6", x"E5E4E3E2",
									 -- x"E4E7E8E8", x"E9EBECEB", x"EEF2F4F6", x"FBFCFBFE", x"FDFDFCFA", x"F9F9F8F8", x"F6F7F7F5", x"F3F2F1F2",
									 -- x"EEEEEDED", x"ECECEAE9", x"EAE9E7E5", x"E3E1DFDE", x"D9D7D4D2", x"D0CFCECD", x"CAC7C5C4", x"C3C2C3C6",
									 -- x"C2C2C4C3", x"BFC1C2BF", x"C0BDBDBD", x"BCB8B6B5", x"BAB7B3B0", x"ADABA8A6", x"A9A7A3A0", x"9E9D9A97",
									 -- x"90929390", x"8D8B8987", x"85807D7C", x"79797772", x"6E6B6966", x"635E5C5B", x"595A5A59", x"5D626260",
									 -- x"60666663", x"65696D70", x"6E717476", x"787A7977", x"7E7E7D7D", x"7C7D7F80", x"7E7C7D7D", x"78767673",
									 -- x"6E6F6E6D", x"6E71706E", x"70707273", x"72707073", x"6F707170", x"6F6E6F70", x"76717175", x"7573757B",
									 -- x"7C7A7A7C", x"7D7C7C7D", x"7F7D7D7E", x"81807D7A", x"7F7C7D82", x"83818285", x"81858B90", x"9396999A",
									 -- x"97999A99", x"999DA2A6", x"A6A5A8B0", x"BAC2C9CD", x"D2CECCCC", x"CFCFCBC8", x"C2C2BFB9", x"B6B6B5B4",
									 -- x"B3AFADA8", x"A19F9C96", x"93959593", x"908F8C8A", x"87858382", x"85878480", x"7C7B7873", x"706D6863",
									 -- x"66666564", x"65676663", x"65646261", x"605E5B58", x"5A595A5A", x"59565556", x"55555554", x"54535251",
									 -- x"CFCFCFCD", x"C9C4C0BE", x"B6B5B4B3", x"B2B1AFAE", x"A8A8A6A5", x"A4A3A2A2", x"A2A5A6A4", x"A4A7A7A4",
									 -- x"A6A7A9AA", x"ABACADAE", x"B3B7B7B6", x"B5B1ACAD", x"AAABADAE", x"ADACA9A8", x"A9ACAFB0", x"B0AFADA9",
									 -- x"AEACA9A8", x"A8A7A4A1", x"A2A4A3A0", x"9FA09F9C", x"97979693", x"9393918D", x"8A8A867F", x"7A79797A",
									 -- x"78746F6C", x"6B6B6B6A", x"69696969", x"69696969", x"68686868", x"68686868", x"67676869", x"69686767",
									 -- x"66646364", x"65625F5E", x"5D5D5D5C", x"5A595B5D", x"5A5C5B5A", x"5B5E5F5E", x"61615F5D", x"5E62625E",
									 -- x"65656669", x"6C6E6E6E", x"716D6968", x"68696968", x"676B6E6D", x"6C6D7071", x"6F757978", x"7B80817E",
									 -- x"807E8085", x"84808288", x"85888D91", x"93949596", x"9DA0A0A1", x"A6A7A7AA", x"AAABACAE", x"AFB0B0B0",
									 -- x"B2B3B3B3", x"B4B8BEC3", x"C2C3C6CA", x"CED2D6D8", x"D9D9D8D7", x"D7D7D7D7", x"D7DADEE0", x"E0DFDFDE",
									 -- x"D9DBD7D1", x"D1D2D3D7", x"DADDE0E0", x"DDDBDCDE", x"DFDDD9D6", x"D5D7DBDE", x"E0E2E5E8", x"E9EBEDEF",
									 -- x"F1F0EEED", x"ECECEDED", x"EDEEEDE9", x"E8E9ECED", x"EEEDEBE8", x"E5E6E8EB", x"E9EAEBEA", x"E9E7E5E3",
									 -- x"E3E5E6E5", x"E6E9EBEB", x"EEF0F0F3", x"FAFCFBFD", x"FDFCFBFA", x"F9F8F7F7", x"F7F7F7F5", x"F2F0EFEF",
									 -- x"ECECEBEB", x"EBEAE9E8", x"E7E6E5E3", x"E1DFDDDD", x"D8D6D3D0", x"CECDCBCB", x"C8C5C3C2", x"C2C1C1C3",
									 -- x"C0C0C1BF", x"BBBCBDB9", x"BCBABABB", x"BAB5B2B2", x"B4B1AEAD", x"ADAAA6A2", x"A6A5A19D", x"9B9B9893",
									 -- x"8D91928E", x"8A888684", x"84807F7D", x"76737473", x"716B6764", x"5F5A5A5D", x"5656575B", x"61666767",
									 -- x"646B6962", x"62666A6E", x"73747373", x"74767572", x"74797F82", x"82818080", x"807D7D7C", x"78767672",
									 -- x"706F6E6E", x"71757470", x"71707273", x"716E6F72", x"6E6F6F6E", x"6D6E7275", x"726F7177", x"78737378",
									 -- x"7C797777", x"78777676", x"79777778", x"7A7A7978", x"7B7A7B7E", x"807F7F7F", x"83888E94", x"9A9FA3A5",
									 -- x"A3A7A6A1", x"9DA0A6AA", x"AAA7A9B5", x"C0C8D0D6", x"D6D4D2D2", x"D1D0CECD", x"CFCFCAC3", x"BEBCBBB9",
									 -- x"B9B3AFA9", x"A4A2A099", x"979C9D98", x"92908F8C", x"8C898686", x"898B8883", x"80807E79", x"75726D68",
									 -- x"696A6A68", x"68696866", x"69666565", x"6564605C", x"5C5C5E60", x"5E5A5857", x"56575757", x"57575655",
									 -- x"CCCCCBCA", x"C7C3BFBC", x"BCB8B3B1", x"B2B1AEAA", x"A6A6A6A7", x"A6A3A2A2", x"A0A2A4A3", x"A1A1A3A6",
									 -- x"A2A5A5A4", x"A4A7A9A9", x"A9ABAEB0", x"AFADADAD", x"ABA9A7A8", x"AAABA9A7", x"A7ACB0AE", x"ADAEACA9",
									 -- x"AEADABA9", x"A9A8A7A5", x"A3A3A3A1", x"A0A09E9B", x"9E9C9A97", x"93909193", x"8C8C8980", x"78767677",
									 -- x"776E6C6E", x"6E6D6C69", x"6866696E", x"6C6A6A67", x"69686767", x"68686868", x"6B696767", x"68696867",
									 -- x"69686563", x"61605F5F", x"5C5E5F5E", x"5B595A5C", x"5B5B5C5C", x"5D5E5F5F", x"5E5E6061", x"62636669",
									 -- x"66696B6E", x"73777875", x"7975706F", x"6E6D6D6D", x"6D727574", x"72737576", x"75787B7D", x"7E808386",
									 -- x"87848488", x"8A898A8D", x"8B8E9194", x"9597999B", x"A0A4A5A5", x"A9B0B3B3", x"B1B0B1B2", x"B3B3B6BA",
									 -- x"B9BAB7B7", x"BDC0C0C3", x"C5C6C9CF", x"D4D6D9DC", x"DDDBD8D8", x"DADBDBDA", x"D9DEE1E1", x"E1E2E2E0",
									 -- x"DCDAD7D2", x"CFD0D4D7", x"DDE0DEDC", x"DDDCDCE0", x"DFDAD8DB", x"DCDADADD", x"E0E5E8EB", x"EFEEECEE",
									 -- x"F1F1F0EF", x"EDEBEAEA", x"EBEDEDEB", x"E9E9EEF2", x"F3EEEBE9", x"E6E3E6EC", x"EEEEEEEE", x"ECEAE7E4",
									 -- x"E4E7E8E7", x"E5E5E9EC", x"ECEEF1F5", x"F8FBFCFD", x"FDFBF9F9", x"F8F6F7F9", x"F6F5F4F3", x"F2F1EEED",
									 -- x"EDECEBEA", x"E9E8E8E8", x"E4E3E2E1", x"E0DEDBD9", x"D6D3D0CF", x"CFCEC9C5", x"C5C5C4C1", x"C0C1C1C0",
									 -- x"C0BEBDBC", x"BBB9BBBF", x"BAB9B9B9", x"B8B4B1B2", x"B3B2AAB0", x"B0A9AAA3", x"A9A1A19E", x"96999B90",
									 -- x"86888F89", x"84888684", x"83827F79", x"726E7072", x"73696161", x"5F5A5B61", x"58525259", x"5E5E6267",
									 -- x"63636260", x"6165696A", x"6C72716F", x"74747173", x"78818688", x"867F7A7B", x"78777777", x"75727171",
									 -- x"6D6C6C6F", x"72747270", x"6F6D736E", x"6A6A656B", x"70706C71", x"6F747173", x"7674766F", x"726E7474",
									 -- x"77797A78", x"7675736F", x"74727274", x"7372767B", x"75737579", x"7C7C7F84", x"898F9598", x"9A9FA3A5",
									 -- x"A5AFABA5", x"AAABAAAF", x"AEACADB7", x"C4CACED6", x"D9D5D2D3", x"D3D1D1D3", x"D1D1CEC9", x"C8C9C4BE",
									 -- x"BDBAB5B1", x"ADA9A5A2", x"A0A09B97", x"97999792", x"92929291", x"908F8C8B", x"8984807D", x"79757170",
									 -- x"70706F6D", x"6C6E6F6F", x"6E6B696A", x"6A676361", x"61666661", x"60625F58", x"5D5B5959", x"5B5C5A57",
									 -- x"CAC9C7C6", x"C4C1BEBC", x"BCB8B3B1", x"B0AFABA8", x"A8A5A3A3", x"A29F9E9F", x"9FA0A1A1", x"A0A0A1A2",
									 -- x"A2A3A2A0", x"A1A4A5A4", x"A5A7A9AB", x"ABABABAB", x"A8A7A6A6", x"A7A8A8A8", x"A5A8ABAB", x"ABABABAA",
									 -- x"ADACAAA9", x"A9A8A8A7", x"A4A1A1A3", x"A29E9C9D", x"99979594", x"92919194", x"8F8F8C85", x"807D7B79",
									 -- x"79747373", x"6F6E6E6C", x"6C68696C", x"6B6A6B69", x"68676666", x"6769696A", x"6A696869", x"6B6B6A69",
									 -- x"68676563", x"61605F5E", x"5E5F605E", x"5C5A5B5D", x"5A5A5A5A", x"5A5C5D5E", x"5F616363", x"63646768",
									 -- x"676B6F72", x"767A7D7D", x"78757578", x"7B7A7775", x"767A7C7D", x"7C7D7D7B", x"7A7D7F81", x"8284878A",
									 -- x"8C8A8A8D", x"8F909193", x"93959799", x"9B9DA0A2", x"A6AAACAC", x"B0B7BAB9", x"B8B8BABC", x"BDBCBEC1",
									 -- x"C0C0BCBB", x"C0C2C3C5", x"C9CACDD2", x"D5D8DCE1", x"E0DDDAD9", x"DADBDCDD", x"DEE2E4E3", x"E3E4E4E3",
									 -- x"DEDCD7D2", x"CFCFD2D5", x"DBDFDEDD", x"DEDDDCDF", x"DDDAD9DB", x"DCDBDDE1", x"E4E9EBED", x"F1F1EFF1",
									 -- x"F0F0F0EF", x"EEECECEB", x"ECEDEDEB", x"E9EAEDF0", x"F2EDE9E9", x"E9E8EAEE", x"F0F0EFEE", x"EDEBE9E7",
									 -- x"E6E7E8E7", x"E5E6E8EB", x"ECEEF1F4", x"F7F9FAFB", x"FDFAF9F9", x"F7F5F5F7", x"F5F4F3F2", x"F0EEECEB",
									 -- x"EBEAE9E8", x"E7E7E7E7", x"E4E2E0DF", x"DDDBD8D6", x"D3D0CECD", x"CFCFCCC9", x"C4C4C3C1", x"C0C1C1BF",
									 -- x"BEBCBCBC", x"B9B6B6B7", x"B6B5B6B8", x"B7B4B0AF", x"B1B1AAAD", x"ADA7A9A5", x"A5A2A3A1", x"99999993",
									 -- x"89878C87", x"81838281", x"83827F7B", x"75716F6F", x"6E696361", x"5F5C5B5C", x"5953535A", x"5D5B5A5D",
									 -- x"5D5B5C60", x"64646466", x"6A6D6D6F", x"75797B7D", x"808B8E89", x"85817C7B", x"75747576", x"75716F6F",
									 -- x"6B6B6B6D", x"7071706F", x"726E736E", x"6C6E686C", x"6B6D6C72", x"70736E6F", x"70727375", x"74747170",
									 -- x"75767675", x"74757370", x"71727170", x"6F707171", x"77747477", x"797A8087", x"8B8F9398", x"9DA3A7A8",
									 -- x"B0B0B0AD", x"ACAFAFAA", x"AAACB0B8", x"C2C6CDD8", x"D6D5D5D5", x"D4D2D3D5", x"D3D4D2CD", x"CCCDC9C3",
									 -- x"C4C0BCB9", x"B6B0A8A1", x"A3A2A0A0", x"A2A29E99", x"9A999999", x"99989694", x"8D898481", x"7C767270",
									 -- x"7272716E", x"6D6E6F6E", x"6F6C6A6C", x"6D6C6967", x"696A6A69", x"68666461", x"605E5B5B", x"5D5E5C5A",
									 -- x"C5C3C1C0", x"C0BFBDBC", x"BAB8B4B1", x"AEABA8A6", x"A9A5A2A1", x"A09F9E9F", x"9D9D9D9D", x"9D9D9D9E",
									 -- x"A2A2A09F", x"9FA1A1A1", x"A4A3A4A5", x"A6A6A6A5", x"A4A5A5A4", x"A4A5A8AA", x"A5A5A5A7", x"A7A7A8AB",
									 -- x"AAA8A7A6", x"A6A7A7A7", x"A7A1A1A4", x"A49E9C9F", x"95939192", x"92919193", x"90908E8A", x"8784807D",
									 -- x"7B7A7A77", x"71707270", x"706B6A6C", x"6A6B6D6B", x"6A696867", x"686A6B6B", x"6A6A6A6C", x"6E6E6D6C",
									 -- x"68676563", x"62605F5E", x"5D5D5E5C", x"5A5A5A5B", x"5B5A5958", x"595B5D5F", x"61646664", x"64676868",
									 -- x"6B70767A", x"7D818587", x"827D7A7D", x"82848383", x"82838484", x"85868583", x"80828485", x"86888C8E",
									 -- x"90919292", x"94979898", x"9B9C9EA0", x"A2A5A8AA", x"ACB0B3B4", x"B8BDC0BF", x"BFBFC2C5", x"C5C4C5C6",
									 -- x"C5C6C2C0", x"C4C6C6CA", x"CFD0D3D6", x"D8DAE0E5", x"E4E1DEDC", x"DBDCDEE0", x"E1E3E4E3", x"E2E3E3E3",
									 -- x"E1DDD8D2", x"CFCFD0D2", x"DADDDEDD", x"DEDCDBDD", x"DCDADADC", x"DCDCDFE4", x"E9EDEEEF", x"F1F1EFF1",
									 -- x"EFEEEEEE", x"EDEDECEC", x"EDEDECEB", x"EBEBEDEE", x"F2EDE9EA", x"ECECEDF0", x"F1F0EFEE", x"EEEDECEB",
									 -- x"E8E8E8E7", x"E6E6E7E8", x"ECEDEFF2", x"F5F7F8F8", x"FAF8F7F7", x"F6F5F4F5", x"F4F2F1F0", x"EEECEAE9",
									 -- x"EAE9E8E7", x"E6E5E5E6", x"E2E0DDDB", x"D9D7D5D4", x"D3D0CCCC", x"CCCCC9C6", x"C5C5C4C1", x"C0C0BFBE",
									 -- x"BBBBBBBB", x"B8B4B2B2", x"B4B2B2B4", x"B5B4B1B0", x"B0B1ADAF", x"AFAAAAA7", x"A0A3A5A1", x"9A969391",
									 -- x"89828581", x"7C7D7B7D", x"807D7A76", x"73706D6B", x"6B68635E", x"5C5C5B5A", x"5B56555A", x"5D5A5959",
									 -- x"5853545B", x"605F5F62", x"68696E73", x"79828888", x"89949488", x"827F7A76", x"72717273", x"726F6D6D",
									 -- x"6F6F6E6E", x"6D6D6D6C", x"716E706E", x"6E706B6B", x"6B6D6A6E", x"6B717275", x"70716D74", x"71797678",
									 -- x"73737271", x"7273726F", x"70716F6B", x"6B6F706D", x"7675777A", x"7C7F878F", x"9396999F", x"A5ABADAB",
									 -- x"B0ADB2B2", x"ABB0B5AC", x"ABB2B7BD", x"C2C5CEDB", x"D8DBDCDA", x"D8D7D7D6", x"D5D8D7D4", x"D2D2CFCB",
									 -- x"C6C3C0C0", x"C0BCB4AC", x"AAA6A4A7", x"A9A8A4A1", x"A2A1A1A2", x"A3A2A09D", x"938E8A87", x"827B7673",
									 -- x"75767472", x"71717170", x"706D6C6E", x"70706F6E", x"706C6B6D", x"6C686668", x"66635F5F", x"5F605F5E",
									 -- x"BEBEBEBD", x"BCBBBCBC", x"B9B7B4B0", x"ADA9A7A5", x"A7A3A1A1", x"A1A0A0A0", x"9A999899", x"9A9B9A9A",
									 -- x"A0A2A2A2", x"A0A0A1A1", x"A5A3A1A1", x"A1A09F9E", x"9F9F9FA0", x"A0A2A4A6", x"A5A2A2A4", x"A5A3A4A8",
									 -- x"A5A4A2A2", x"A2A4A5A6", x"A6A2A1A2", x"A19D9B9C", x"97949292", x"93919090", x"8E8E8D8B", x"88868482",
									 -- x"7E7F7F7A", x"74757874", x"756F6D6D", x"6B6C6E6B", x"6D6C6B6A", x"6A6B6B6B", x"6C6C6C6D", x"6F706F6F",
									 -- x"6A686765", x"63616060", x"5D5D5C5B", x"5A5A5A5A", x"5C5B5A5A", x"5B5D5F60", x"61656765", x"65686968",
									 -- x"6D72797F", x"83878B8D", x"8E898687", x"8A8B8B8C", x"8F8E8D8C", x"8B8C8D8D", x"8888898A", x"8B8E9194",
									 -- x"969A9B99", x"9A9EA09F", x"A2A4A7AA", x"ACAEB0B1", x"B1B5B8BB", x"BFC3C5C4", x"C5C5C7CA", x"CBCACACB",
									 -- x"CBCCC9C7", x"CACCCDD1", x"D5D7DADB", x"DCDEE2E6", x"E8E6E3E0", x"DEDEE0E1", x"E2E3E3E3", x"E2E2E1E0",
									 -- x"E3DFD9D3", x"D0CFCFD0", x"D9DDDDDC", x"DCDAD8DA", x"DCDBDCDC", x"DBDBDFE4", x"ECEFEEED", x"EFEDEBED",
									 -- x"ECECECEC", x"ECEDEDEC", x"EDECEBEB", x"ECECEDEC", x"F2EEEBEB", x"ECECEDEF", x"EFEFEEEE", x"EEEFEEED",
									 -- x"EAE9E8E7", x"E7E7E7E6", x"EBECEEF1", x"F3F5F6F7", x"F7F6F6F6", x"F5F4F4F4", x"F2F1EFEE", x"EDEBEAE8",
									 -- x"E9E8E7E6", x"E5E5E5E5", x"DFDDDAD7", x"D5D4D3D3", x"D2D0CECD", x"CDCCC9C6", x"C7C6C5C2", x"BFBEBCBB",
									 -- x"BBBABAB8", x"B6B4B2B1", x"B4B1AEAF", x"B2B3B2B1", x"AEAFAEB1", x"B1AEAAA7", x"A0A5A49F", x"99928D8D",
									 -- x"887E7F7E", x"7A78777A", x"7D797470", x"6D6C6C6B", x"6B655F5A", x"5958595A", x"5C575557", x"5A5B5B5C",
									 -- x"57535155", x"595B5F63", x"67676F77", x"7B86908E", x"92989388", x"827E7773", x"73717070", x"6F6D6C6D",
									 -- x"6F6F6E6D", x"6B6A6B6C", x"6B6B6D6C", x"6D6E6B69", x"6D706C6E", x"6A717277", x"73716C70", x"70777779",
									 -- x"77757271", x"7172706F", x"6F6F6C6A", x"6B6E7273", x"73767C82", x"85899098", x"9DA0A5A9", x"ADB0AFAD",
									 -- x"A9AAADAB", x"A4A8AFAE", x"B1BAC1C4", x"C7CAD3DF", x"E0E4E5E2", x"DFDFDCD8", x"D8DBDCDA", x"D7D7D5D3",
									 -- x"CBC7C3C2", x"C3C2BEBA", x"B4ABA6A7", x"AAA9A7A6", x"A6A5A5A7", x"A9A9A6A3", x"99938E8C", x"89837D78",
									 -- x"79797876", x"76777675", x"75737173", x"75757575", x"74716E6E", x"6E6B696A", x"6A666362", x"62616162",
									 -- x"B9BBBCBB", x"B8B6B6B8", x"B5B5B3AF", x"ACA8A6A5", x"A2A09FA1", x"A19F9D9C", x"97969495", x"97989797",
									 -- x"9C9FA3A3", x"A19E9FA1", x"A5A2A09E", x"9D9C9A98", x"97969798", x"9A9B9C9C", x"A19F9FA2", x"A3A1A0A3",
									 -- x"A0A09F9E", x"9FA0A2A3", x"A1A2A19E", x"9D9E9C99", x"97949293", x"93918F8F", x"8B8C8C89", x"86848689",
									 -- x"8785837E", x"797C7D78", x"78737271", x"6F70706B", x"6D6C6B6B", x"6B6B6B6A", x"6D6D6D6D", x"6E6F6F70",
									 -- x"6C6B6866", x"64636363", x"605F5E5D", x"5D5C5C5C", x"5C5C5C5C", x"5D5E5F60", x"60646665", x"65686A69",
									 -- x"6D717880", x"868A8D8F", x"91929597", x"96939191", x"999B9C9A", x"97959698", x"90909091", x"9296999C",
									 -- x"A1A5A6A3", x"A3A6A8A8", x"ABADB2B6", x"B9BAB9B8", x"B9BCBFC3", x"C6C9CACA", x"CDCCCDCF", x"D0CFD0D1",
									 -- x"D0D2D0CE", x"D1D2D4D8", x"D8DBDFE1", x"E2E4E7E9", x"EBEAE8E5", x"E2E1E1E1", x"E3E2E3E3", x"E3E1DFDE",
									 -- x"E2DFDAD4", x"D0CECECF", x"D9DCDBD9", x"D9D6D4D7", x"DADBDDDC", x"DBDBDFE4", x"EAEDECEB", x"ECEBE9EB",
									 -- x"ECEBEBEB", x"EDEEEEEE", x"ECEBEBEB", x"ECEDEDEC", x"EFEDECEB", x"EAEAECEF", x"EEEEEEEE", x"EEEEECEB",
									 -- x"EAE9E7E7", x"E8E7E7E6", x"EAEBEDEF", x"F2F4F6F7", x"F5F6F5F5", x"F4F3F2F1", x"F1F0EEED", x"ECECEAE9",
									 -- x"E7E7E5E4", x"E3E3E3E3", x"DFDDD9D5", x"D2D1D0D1", x"CFCFCFD0", x"D1D0CDCA", x"C8C6C4C1", x"BFBCBBBB",
									 -- x"BDBBB8B5", x"B3B3B2B1", x"B1AFADAD", x"AFB1B0AE", x"ABAAABAD", x"AFB0ACA8", x"A6A6A39E", x"9A938D8E",
									 -- x"8A7E7F7E", x"79767478", x"7A78736F", x"6C6A6969", x"68605A5A", x"59545559", x"59565455", x"56575858",
									 -- x"54565553", x"555D6467", x"67676E74", x"78859293", x"97968F88", x"857F7775", x"7673706F", x"6D6C6C6E",
									 -- x"696A6A69", x"68686A6C", x"64686A6A", x"6A6A6A67", x"6B717175", x"6F726E6D", x"736F706F", x"75747471",
									 -- x"7B787573", x"71706E6D", x"6E6B6B6F", x"6F6E7278", x"767A8086", x"898D949A", x"9EA5ACB0", x"B1B1B1AF",
									 -- x"ADAFA8A1", x"A2A3A5AB", x"B5BFC5C8", x"CDD2DBE4", x"E7E9E9E7", x"E6E6E1DB", x"DBDDDFDD", x"DBD9D9D8",
									 -- x"D6D1CBC7", x"C4C2BFBE", x"BAB1AAAA", x"ABAAA9AA", x"AAA9AAAC", x"AEADAAA7", x"9E97908E", x"8D88817C",
									 -- x"7C7C7B7A", x"7B7C7C7A", x"7D7B7A7B", x"7C7B7A7B", x"7B7A7773", x"7272716D", x"6B676565", x"65656566",
									 -- x"B7B8B9B6", x"B2B0B0B1", x"B1B0AFAC", x"AAA7A5A3", x"A0A0A1A2", x"A09C9998", x"95939191", x"92939494",
									 -- x"95989C9E", x"9C999A9C", x"9E9E9C9B", x"9A989695", x"93929293", x"95969594", x"9A999B9D", x"9F9E9D9D",
									 -- x"9C9C9C9C", x"9C9D9EA0", x"9EA2A19C", x"9C9F9F99", x"95939293", x"92908E8E", x"8C8C8C8B", x"8786898D",
									 -- x"8F8B8885", x"8282827C", x"7B777777", x"7576736D", x"6C6B6A6A", x"6A6B6B6A", x"6D6C6C6C", x"6C6D6E6F",
									 -- x"6D6C6967", x"65646363", x"615F5D5C", x"5C5D5C5B", x"5B5B5C5D", x"5E5F5F5F", x"60626465", x"6667696B",
									 -- x"6F727880", x"888D9194", x"9597999A", x"9896989B", x"9FA2A6A7", x"A39E9D9E", x"98979696", x"999DA1A4",
									 -- x"A9ADAEAD", x"ABACAFB1", x"B2B5BABF", x"C2C3C1BF", x"BFC1C5C8", x"CCCECFCE", x"D2D0D0D1", x"D3D3D3D5",
									 -- x"D4D7D5D3", x"D4D5D6DC", x"DCDFE3E6", x"E9ECEDEC", x"EEEDECEA", x"E8E6E4E3", x"E3E1E1E2", x"E1DEDBDA",
									 -- x"DEDDD9D5", x"D0CECECF", x"D7DAD9D8", x"D8D5D3D5", x"D9DBDDDD", x"DCDDE0E4", x"E6E9E9E9", x"ECEBEAEC",
									 -- x"ECEBEAEB", x"EEEFF0EF", x"EDECEBEB", x"ECECECEC", x"EBEBEBEA", x"E9E9ECEE", x"EFEEEEED", x"EDEBE9E7",
									 -- x"E9E8E8E8", x"E8E8E7E6", x"E9EAECEE", x"F0F3F4F5", x"F5F6F6F4", x"F3F2F0ED", x"EFEEEDEC", x"EBEBEAE9",
									 -- x"E5E4E3E2", x"E1E0E0E0", x"DFDDD9D4", x"D0CECECE", x"CFCFD0D1", x"D0CECAC6", x"C5C3C1BF", x"BEBCBBBC",
									 -- x"BDBBB7B3", x"B1B1B1B0", x"ADADACAC", x"ADADAAA6", x"AAA8ABA9", x"ACB2AFAF", x"ABA7A3A0", x"9B979594",
									 -- x"8A80807C", x"75727074", x"76757370", x"6C686462", x"635B585C", x"5B535155", x"55565756", x"55545250",
									 -- x"4C535654", x"565E6464", x"67696C6F", x"73809198", x"96928A85", x"837D7676", x"77747271", x"6F6D6D6E",
									 -- x"6B6B6B69", x"66656667", x"5F666567", x"67676A66", x"686E6E72", x"6F74706F", x"726E716E", x"79787E7B",
									 -- x"7D7A7674", x"706D6C6D", x"6F6B6E76", x"77727278", x"7E818486", x"898D9398", x"9DA7B0B3", x"B2B2B3B4",
									 -- x"B6B4A7A1", x"ACAFACB2", x"B8C2C7CA", x"D2D9E0E7", x"E8E7E7E8", x"EAEAE5E0", x"DEDFDFDE", x"DCDBDBDB",
									 -- x"DBD7D1CC", x"C7C3C0BE", x"BDB8B2B1", x"B1B0AEAD", x"AEAFB0B2", x"B2B0AEAC", x"A29B9490", x"8E898480",
									 -- x"8281807E", x"7F81817F", x"807F7F81", x"82807F80", x"82817D78", x"78797772", x"6C69686A", x"6B6A6A6C",
									 -- x"B4B3B1AF", x"ADADACAC", x"ADACAAA8", x"A7A4A2A0", x"9E9FA1A2", x"9E989595", x"94928F8D", x"8D8E8F90",
									 -- x"8F8F9194", x"95939395", x"96979898", x"96949392", x"92929291", x"91919192", x"93959696", x"98989794",
									 -- x"98989998", x"9798999B", x"9C9D9C99", x"989A9996", x"93929393", x"928F8F90", x"8E8D8E8E", x"8C8A8A8D",
									 -- x"908B8B8C", x"89878581", x"7D7B7B7C", x"7B7C7971", x"6E6C6A69", x"696B6C6C", x"6A6A6B6B", x"6B6B6C6C",
									 -- x"6B6A6968", x"66646261", x"605D5A5A", x"5B5C5B5A", x"5B5C5D5E", x"5F5F5F5F", x"62616366", x"6766686D",
									 -- x"6E71777F", x"868C949A", x"9F9D9B9A", x"999A9FA4", x"A4A6AAAC", x"AAA5A3A3", x"A19F9E9E", x"A1A6AAAD",
									 -- x"B0B2B4B5", x"B3B1B5B9", x"BABCBFC4", x"C7C9C8C7", x"C6C8CBCE", x"D1D2D3D3", x"D4D2D2D3", x"D5D5D5D5",
									 -- x"D5D9D9D8", x"D9D9DBE0", x"E2E5E8EB", x"EFF2F2F0", x"F1EFEEED", x"ECEBE8E7", x"E5E2E0E0", x"DFDBD8D7",
									 -- x"D8D9D8D5", x"CFCDCED0", x"D3D7D8D7", x"D8D6D3D5", x"DBDCDEDE", x"DDDEE0E2", x"E2E6E7E8", x"EBEBEAEC",
									 -- x"ECEAE9EA", x"EDEFF0EF", x"EEEDEDEB", x"EBEAEBEB", x"E9EAE9E9", x"E9EAECEC", x"EFEEEDEB", x"EBE9E8E7",
									 -- x"E7E8E8E8", x"E8E8E8E8", x"E9E9EAEC", x"EEF0F2F3", x"F3F5F5F4", x"F2F2F0ED", x"EEECEBEA", x"E9E8E8E7",
									 -- x"E3E3E1E0", x"DFDFDFDF", x"DCDBD8D3", x"CFCDCDCE", x"D3D2D1D0", x"CECAC5C1", x"C3C0BEBD", x"BBB9BABC",
									 -- x"BBBAB7B4", x"B3B3B1AE", x"ADAEADAA", x"A9A9A7A4", x"A7A8AFAC", x"ACB1ADB0", x"ADA4A3A1", x"9A989A97",
									 -- x"8B83827B", x"72707074", x"74716F6E", x"6C69635F", x"5F5B595B", x"5A555252", x"51555653", x"504F4E4D",
									 -- x"4B515657", x"5A5E605F", x"62686A69", x"6F7A8996", x"96958C81", x"7D797574", x"74737475", x"736F6D6C",
									 -- x"6F6E6C69", x"66646463", x"5E635F61", x"63656A65", x"666A696D", x"6D767575", x"6D6C6D71", x"7A81888A",
									 -- x"817F7D7A", x"76727275", x"7873747B", x"7F7D7A7B", x"8386888A", x"8D919598", x"9FA8B0B1", x"B0B0B2B4",
									 -- x"B5B0AAAB", x"B2B8BBBE", x"C2CCCFD0", x"D6DDE2E6", x"E6E5E5E8", x"EBE9E7E5", x"E0E0DFDE", x"DDDBDBDB",
									 -- x"DBD6CFCB", x"C8C7C4C2", x"BFBDBAB6", x"B4B3B1AF", x"B0B2B4B5", x"B4B1AFAE", x"A39F9994", x"8F8A888A",
									 -- x"8A898784", x"85878684", x"82828488", x"89888787", x"87827E7D", x"7C7B7876", x"716F6F71", x"716E6D70",
									 -- x"B1ADA9A8", x"AAACACAA", x"AAA9A6A5", x"A4A29F9C", x"999B9E9F", x"9A949192", x"93918E8B", x"8A8B8C8E",
									 -- x"8D8A898D", x"90908F8F", x"90929595", x"93919090", x"9091918F", x"8C8B8E91", x"90929391", x"9294918D",
									 -- x"94959595", x"94949596", x"98969493", x"928F8E8E", x"93939495", x"93908F91", x"8F8E8F91", x"918D8B8B",
									 -- x"8C888C90", x"8D898785", x"7F7D7E7F", x"7F807D75", x"73706C69", x"696B6D6E", x"67686A6A", x"6A6A6A6B",
									 -- x"68696968", x"6663615F", x"615E5B5A", x"5C5D5C5A", x"5D5D5D5E", x"5F606061", x"64616267", x"6765686E",
									 -- x"6A6E747B", x"8187929D", x"A6A4A2A2", x"A1A1A3A6", x"ABA9AAAC", x"ACAAA9AA", x"AAA8A6A7", x"AAAFB4B7",
									 -- x"B7B7BABC", x"BAB7BBC1", x"C2C3C4C8", x"CBCECFCF", x"CDCED1D5", x"D7D8D9D9", x"D7D5D4D6", x"D8D7D7D7",
									 -- x"D8DDDEDE", x"DFE0E2E8", x"E9EBECEE", x"F2F5F4F1", x"F3F1EEEE", x"EFEEECEA", x"EAE6E2E1", x"DFDBD8D8",
									 -- x"D4D6D7D4", x"CFCCCDD0", x"CFD5D7D8", x"DAD8D5D6", x"DDDFE0DF", x"DEDEDFE0", x"E1E5E5E6", x"EAE9E8EB",
									 -- x"EAE8E7E8", x"EBEEEEEE", x"EFEFEEEC", x"EAE9E9EA", x"EBEAE8E8", x"E9EBEBEA", x"EFEDEBEA", x"E9E9E9E9",
									 -- x"E6E7E8E8", x"E8E8E8E9", x"E8E9EAEB", x"EDEFF0F1", x"F1F3F4F3", x"F3F3F1EE", x"EDEBE9E8", x"E7E6E6E5",
									 -- x"E4E3E2E1", x"E0DFDFDF", x"D9D8D5D2", x"CFCDCECF", x"D5D4D3D2", x"CFCCC8C5", x"C3BFBCBB", x"B9B7B8BA",
									 -- x"B8B9B8B6", x"B6B6B3AF", x"B2B1ADA7", x"A5A6A7A6", x"A3A7B4AF", x"ABADA7AB", x"ABA1A2A1", x"97959A97",
									 -- x"8E87867C", x"73737579", x"76716D6C", x"6E6D6863", x"5F5D5A58", x"57565452", x"4B50514D", x"494A4D4D",
									 -- x"5253575C", x"5F5E5E5E", x"59646665", x"6B727E8D", x"999C9281", x"79787573", x"71727578", x"77716C6A",
									 -- x"6A696866", x"66656464", x"5D61595C", x"60636A63", x"646B6B71", x"70787370", x"64696C79", x"7C868588",
									 -- x"88878685", x"807C7E81", x"827D797C", x"83878581", x"83878C91", x"95989A9A", x"A1A8ADAD", x"AAAAACAE",
									 -- x"ADA9AFB2", x"AEB4C0C1", x"CED7D9D6", x"D9DDE0E3", x"E6E4E5E9", x"EAE8E7E9", x"E2E0DFDE", x"DDDCDBDB",
									 -- x"DCD4CBC7", x"C7C7C6C3", x"C1C1BDB5", x"B2B2B2AF", x"B0B3B5B5", x"B3B0AEAE", x"A2A19E98", x"908B8E93",
									 -- x"92908D8A", x"8A8B8A88", x"85868A8F", x"92919090", x"8A827E81", x"817B787A", x"77757577", x"76716E70",
									 -- x"ACA9A7A7", x"A5A2A4AA", x"A7A5A3A0", x"9E9C9A98", x"92949698", x"96918F8F", x"908C8989", x"8A898888",
									 -- x"8B87888A", x"888B9193", x"93939292", x"9190908F", x"9090908E", x"8C8C8C8D", x"8F8D8C8E", x"8D8B8C90",
									 -- x"90908F8E", x"8E8E8F8F", x"8F8E8F91", x"92908F8F", x"90929392", x"908F9092", x"928F8F92", x"93908E8E",
									 -- x"8D909291", x"8F8E8C8A", x"87807D80", x"807C7B7E", x"78726D6D", x"6F6F6E6D", x"6C686565", x"66656667",
									 -- x"6B696766", x"64616163", x"625D5A5B", x"5D5E5E5E", x"5A5E5E5D", x"5F5E5F64", x"62636567", x"6767696B",
									 -- x"6D727879", x"80898F9C", x"A8A8A8A6", x"A3A4A8AB", x"ABACAEAF", x"AFAFAFB0", x"AEABAFB6", x"B6B1B7C4",
									 -- x"BFBEBEC0", x"C1C1C4C8", x"C3C8CCCF", x"D3D7D5D1", x"D2D1D2D8", x"DCDCDBDB", x"DADADAD9", x"D7D7D8D9",
									 -- x"DBDCDDDE", x"E1E5E9EC", x"EDEDEEEF", x"F1F3F5F7", x"F3F4F4F3", x"F2F2F0EE", x"ECE6E3E4", x"E2DDD9D9",
									 -- x"D2D2D1CF", x"CECFCECB", x"CFD3D6D6", x"D7DADAD8", x"DBDEE2E5", x"E5E4E3E4", x"E4E6E8E9", x"E8E7E7E7",
									 -- x"E6E8E9EA", x"EBEBEDEE", x"EFEDEDEE", x"ECE9E7E7", x"E9E7E6E6", x"E8E9EAE9", x"E8E9EAE9", x"E7E6E7E8",
									 -- x"E6E4E3E3", x"E5E7E8E7", x"E8E8E9EA", x"EBEDEEEF", x"EDEFF1F2", x"F1EFEDEC", x"ECEAE8E7", x"E7E7E6E6",
									 -- x"E3E2E2E2", x"E1E0DFDD", x"DAD5D2D1", x"CECBCDD2", x"D4D2D1D2", x"D7D7D0C8", x"C6C3BFBB", x"BBB9B4AE",
									 -- x"BAB8B8B7", x"B5B0AEAE", x"AEABA5A1", x"A1A3A9AD", x"ACADADAB", x"ABACABA9", x"AEA59C98", x"95918F90",
									 -- x"918B8682", x"7B736E6E", x"6E6F6E69", x"6868645E", x"5B595756", x"5859544E", x"4A4E504D", x"48494D52",
									 -- x"555E6160", x"6364615F", x"635F6969", x"686B7185", x"909A9185", x"78727976", x"746E737A", x"7776736A",
									 -- x"69686969", x"67686660", x"625E5F5E", x"5A606662", x"686A6C6E", x"6E6D6B6A", x"696D6F74", x"7D828488",
									 -- x"8F8D8A86", x"817E7F81", x"84828081", x"83868888", x"8E919096", x"97949CA0", x"A2AAABA9", x"ABACABAB",
									 -- x"ADACB2B9", x"B7B9C5D1", x"D7DADCDB", x"D7D7DBE0", x"E3E4E7EA", x"EAE8E6E4", x"DDDDDDDD", x"DDDCD8D5",
									 -- x"D4D1CDC9", x"C7C6C6C7", x"C2C0BBB4", x"B2B8B7AD", x"B6B4B5B6", x"B2B0ADA7", x"A29F9D9A", x"94949898",
									 -- x"93959391", x"92949089", x"8A8C8F91", x"93928F8A", x"89888683", x"807F7E7C", x"7F7C7977", x"77787776",
									 -- x"A7A6A6A7", x"A4A0A0A4", x"A2A19F9D", x"9B989593", x"908E8E8F", x"8E8C8A8A", x"8A878687", x"88878686",
									 -- x"8582868A", x"898B8F90", x"8F8F9091", x"91919191", x"8F8F8F8E", x"8C8C8C8D", x"8C8A898D", x"8D8B898B",
									 -- x"8C8B8C8C", x"8C8D8D8E", x"8E8D8D8E", x"8E8D8C8E", x"9090908E", x"8B8B8C8E", x"92909091", x"91908F90",
									 -- x"91949694", x"92908D8B", x"8A848080", x"7F7D7C7E", x"7A746F6F", x"706F6D6C", x"6C686565", x"67666666",
									 -- x"68666666", x"64616162", x"645F5C5B", x"5D5D5D5E", x"5B5F5F5E", x"5F5E5E63", x"63636465", x"6565686B",
									 -- x"70727777", x"7F898F9B", x"A4A6A7A6", x"A3A3A6A9", x"ACAEB1B5", x"B8B9B9B9", x"B7B8BABB", x"BAB9BDC2",
									 -- x"C6C4C3C4", x"C4C5C8CC", x"CCCDCED0", x"D4D8DAD9", x"DAD8D9DD", x"E0DFDEDE", x"DFDEDCDB", x"DBDCDBDB",
									 -- x"D8D9DCDF", x"E3E7EBED", x"EEEEEFF1", x"F2F5F7F9", x"F6F6F6F5", x"F5F6F4F2", x"ECE7E4E5", x"E5DFDBDB",
									 -- x"D3D0CDCD", x"CFCFCCCA", x"CED3D7D8", x"DADDDDDC", x"DEE0E3E6", x"E6E6E6E6", x"E5E5E6E7", x"E9E9E8E7",
									 -- x"E6E7E8E9", x"E9EBEEF0", x"EEEDEDEE", x"EDEAE8E9", x"E9E9E9E8", x"E8E8E9E9", x"E7E8E8E7", x"E6E5E6E6",
									 -- x"E5E3E2E2", x"E4E5E6E6", x"E5E6E7E9", x"EBEDEEEF", x"EEEEEEEF", x"F0EFEEEC", x"EDECEAE8", x"E5E4E3E4",
									 -- x"E4E3E2E1", x"E0DFDEDC", x"DAD6D2D1", x"CECCCFD4", x"D6D3D0D0", x"D5D7D4CE", x"CBC9C5C1", x"BEBCB9B5",
									 -- x"B9B6B4B3", x"B2AFADAD", x"ABA7A5A6", x"A4A1A4AB", x"ADACA9A6", x"A5A7A8A7", x"A49F9B98", x"95918F8F",
									 -- x"938D857D", x"77727070", x"6D6E6C67", x"6464625E", x"59595756", x"5757534D", x"4D51514D", x"4B4E5357",
									 -- x"5F646564", x"65625D5C", x"5E5F6968", x"686E707B", x"8A948E84", x"78727773", x"75707379", x"7776736B",
									 -- x"68676867", x"6363635E", x"6261615F", x"5E616260", x"6466686B", x"6C6C6B6A", x"70737579", x"8185868A",
									 -- x"8D898584", x"87898987", x"83858889", x"8A8D9297", x"90989BA0", x"9E9BA3A6", x"A0A4A3A2", x"A8ACAFB3",
									 -- x"B0B4B9BC", x"BCBECAD7", x"D7D8D9D9", x"D9D9DBDD", x"DFE2E5E7", x"E7E5E2E1", x"DBDADADA", x"D9D7D3D0",
									 -- x"D2CDC7C7", x"C9CBC9C6", x"C4C3C1BC", x"B7BABBB4", x"B3B1B3B5", x"B3B1ADA7", x"A7A09C9B", x"9A9B9B97",
									 -- x"9C9D9C99", x"999B9994", x"94949494", x"9494918D", x"8E8D8A87", x"86858585", x"85837F7D", x"7C7C7A78",
									 -- x"A3A2A2A3", x"A19D9C9F", x"9F9F9E9D", x"9A97928F", x"8F8B8888", x"89888788", x"84848587", x"87858485",
									 -- x"82808489", x"88898D8D", x"8D8E8F90", x"91929292", x"8C8C8C8C", x"8B8B8B8C", x"8B878588", x"8A898787",
									 -- x"87878788", x"898A8B8B", x"8D8B8A8B", x"8B8A8A8C", x"8A8A8988", x"88898D90", x"92919090", x"90909192",
									 -- x"94969896", x"94928F8C", x"8C898480", x"7F7F7E7E", x"7B767271", x"71706D6C", x"6B676464", x"65646362",
									 -- x"64646466", x"64626162", x"66615D5C", x"5C5C5C5D", x"5C60605E", x"5F5E5E62", x"64636465", x"6566696D",
									 -- x"71717575", x"7F8A8F9A", x"A2A6AAAA", x"A7A5A6A9", x"ADB0B5BB", x"BFC1C0BE", x"C1C5C6C3", x"C2C6C7C5",
									 -- x"CBCAC9CB", x"CBCBCDD0", x"D4D2D2D4", x"D8DBDFE2", x"E2E1E1E3", x"E5E4E3E3", x"E2E0DDDC", x"DDDDDCDB",
									 -- x"D9DBDEE3", x"E7ECEFF1", x"F0F0F1F1", x"F3F6F9FB", x"F9F9F7F7", x"F8FAF9F6", x"EDE9E7E9", x"E9E4DFDD",
									 -- x"D6CFCBCE", x"D2D1CECC", x"D0D4D8DB", x"DEE0E1E0", x"E1E2E5E7", x"E8E8E7E7", x"E7E6E5E6", x"E8E8E7E6",
									 -- x"E8E8E8E8", x"E9EBEDEF", x"EEEDEDEE", x"EDEBEAEA", x"E7E8E9E9", x"E6E5E5E6", x"E7E6E5E5", x"E5E5E4E4",
									 -- x"E5E3E0E0", x"E1E3E3E3", x"E3E4E6E8", x"EAECEDED", x"EFEDEBEC", x"EEEFEEEC", x"EAEBEBE9", x"E6E5E6E8",
									 -- x"E5E3E1E0", x"DFDDDCDB", x"D9D6D4D3", x"D1CED0D5", x"D6D4D1D2", x"D6D9D7D2", x"CDCCC9C4", x"C1BFBDBB",
									 -- x"B8B4B1B1", x"B0ADABA9", x"ABA5A3A5", x"A29C9EA5", x"ACAAA7A4", x"A2A3A2A1", x"9C9C9B97", x"94928F8C",
									 -- x"8E8C8781", x"7B76716D", x"6B6C6A65", x"62615E5B", x"57575655", x"5554504D", x"5154534E", x"4C52585A",
									 -- x"64666564", x"635D585A", x"5F636B69", x"6A717174", x"87908E88", x"7F787975", x"7270757B", x"7A77736D",
									 -- x"69686966", x"5F5F605D", x"62636160", x"63646262", x"60626568", x"6B6C6D6E", x"7478797D", x"8487878A",
									 -- x"8A8A8989", x"8C8F8C87", x"85898C8E", x"8F92989C", x"929CA0A3", x"A1A0A8AA", x"A8AAA8AA", x"AFB1B2B8",
									 -- x"B5C0C3C2", x"C4C4C9D5", x"D9D7D6D6", x"D8DAD9D8", x"DBDEE1E2", x"E0DEDBDA", x"D5D5D6D6", x"D6D3CFCC",
									 -- x"CBC7C4C5", x"C8CACAC8", x"C4C5C7C5", x"BFBEBEBB", x"B6B2B3B5", x"B4B3B1AB", x"ACA5A1A0", x"9FA1A19D",
									 -- x"A3A5A4A1", x"A0A1A09D", x"9E9D9B98", x"98989693", x"93918E8C", x"8B8A8B8C", x"89868482", x"817F7C7A",
									 -- x"9E9D9D9E", x"9C9A9A9C", x"9C9C9B9A", x"9995918F", x"8C898787", x"87868586", x"81828486", x"86838283",
									 -- x"84818487", x"85878B8B", x"8C8C8D8E", x"8E8E8E8D", x"89898989", x"89898A8A", x"8B868284", x"85848587",
									 -- x"83848485", x"86878888", x"8C8A898A", x"8B8A8B8C", x"89888685", x"868A8F93", x"918F8E8F", x"91939392",
									 -- x"93969797", x"9594928F", x"8C8B8782", x"8081807D", x"7B767373", x"72706D6C", x"68656363", x"62616060",
									 -- x"62626466", x"65626061", x"64615F5E", x"5D5B5B5B", x"5C5F5F5E", x"5F5E5E62", x"63636567", x"68686C70",
									 -- x"6F717576", x"7F898E99", x"A2A8AEAF", x"ABA8A8AA", x"B0B3B7BC", x"C2C4C2BE", x"C6CACCCB", x"CCD0D1CE",
									 -- x"D0D0D2D5", x"D6D5D5D7", x"D9D6D7DB", x"DEDFE3E7", x"E7E6E6E7", x"E8E8E7E7", x"E5E3E1DF", x"DDDCDBDB",
									 -- x"DBDDE1E6", x"EBEFF1F2", x"F2F2F2F2", x"F3F5F8FB", x"FBF9F7F7", x"F9FCFCF9", x"EEECEBEE", x"EEE9E2DE",
									 -- x"D8D0CCD1", x"D5D4D2D3", x"D4D6DADD", x"DFE1E2E2", x"E4E4E6E7", x"E9E9E8E7", x"E9E8E7E6", x"E6E6E6E5",
									 -- x"E9E9E9E9", x"EAEBEDEE", x"F0EFEFEE", x"EDECEAEA", x"E6E7E8E8", x"E6E4E3E3", x"E6E4E3E3", x"E5E6E4E3",
									 -- x"E4E2DFDE", x"DFE0E1E1", x"E2E3E5E8", x"E9EAEAEA", x"EDECEBEB", x"EDEEEEED", x"E9E9E9E8", x"E7E6E7E7",
									 -- x"E5E3E1DF", x"DDDCDAD9", x"D6D5D5D6", x"D3CFCED1", x"D4D4D5D7", x"DBDCD8D3", x"CECDCAC6", x"C5C4C1BF",
									 -- x"B7B3B0B1", x"B0ACA7A5", x"A8A3A09F", x"9E9DA0A5", x"A8A8A8A8", x"A6A4A09E", x"999C9A95", x"908F8C88",
									 -- x"8A8C8A84", x"807C756D", x"6A6A6865", x"63615C56", x"55555452", x"51504F4E", x"5155554F", x"4D52585A",
									 -- x"615F5C5D", x"5D57555B", x"666B706E", x"6F737677", x"7F878B89", x"827C7874", x"71747A7F", x"7C76716E",
									 -- x"69696B68", x"62626666", x"62656160", x"6869666A", x"63646567", x"696B6C6D", x"73777A7E", x"85878587",
									 -- x"868E9393", x"91918E8A", x"8D8C8C8E", x"92959695", x"99A2A3A6", x"A8ACB3B1", x"B2B5B8BC", x"BEB8B6BB",
									 -- x"BECCCDC9", x"CCC9C5CC", x"D9D7D4D3", x"D5D7D6D4", x"D6D9DAD9", x"D6D4D3D2", x"D4D4D4D4", x"D3D0CCC8",
									 -- x"C3C5C6C5", x"C3C4C8CB", x"C8C8CDCE", x"C9C6C6C3", x"C2BBB9B8", x"B7B8B7B3", x"AEABAAA7", x"A2A2A6A6",
									 -- x"A7AAAAA8", x"A6A6A5A4", x"A2A2A09E", x"9E9F9E9B", x"98959392", x"908F8F90", x"8B888686", x"8684807D",
									 -- x"9797999A", x"9A989797", x"95959493", x"92908E8C", x"86868686", x"84818081", x"7D7E8083", x"83818182",
									 -- x"827F8285", x"84848888", x"88888989", x"89888786", x"88888888", x"88898888", x"88848283", x"82808286",
									 -- x"80808183", x"84868788", x"8A89898B", x"8C8B8C8D", x"8B8A8785", x"86888C8F", x"8F8C8B8D", x"92959491",
									 -- x"94969796", x"9594928F", x"8A8B8985", x"8485827D", x"7B777473", x"716E6B69", x"63626363", x"615F5F61",
									 -- x"61626466", x"65615F60", x"605F5F5F", x"5D5B5A5B", x"5C5F5E5D", x"5F5E5E61", x"63646668", x"69696B6E",
									 -- x"6F737979", x"7E868B96", x"A1A7AEB0", x"AEAAA9AA", x"B1B4B8BD", x"C4C8C7C3", x"CACBCED2", x"D5D6D7D8",
									 -- x"D8D8DADE", x"DFE0E2E5", x"E1DFDFE2", x"E3E3E6EB", x"ECEBEAEA", x"EAEAEAE9", x"E9E9E8E5", x"E0DDDDDE",
									 -- x"DCDDE0E5", x"EBF0F2F3", x"F4F5F5F4", x"F3F5F8FB", x"FAF8F6F6", x"F8FCFBF9", x"F0EFEFF2", x"F3EEE5DF",
									 -- x"DAD4D2D5", x"D6D4D5D8", x"D8D9DBDE", x"DFE0E2E3", x"E5E6E8E9", x"EAE9E9E8", x"E9EAE9E7", x"E5E4E6E8",
									 -- x"E9E9EAEB", x"ECEEEFEF", x"F2F2F1EF", x"EDEBEAE9", x"E8E8E8E8", x"E9E8E6E4", x"E5E3E2E3", x"E6E7E5E4",
									 -- x"E3E1DFDE", x"DEDFDFDF", x"E1E3E5E7", x"E8E9E9E8", x"E9EAECEC", x"EBEBECED", x"EBE9E6E5", x"E6E5E3E1",
									 -- x"E5E3E0DE", x"DDDBDAD9", x"D5D3D2D3", x"CFCBCACD", x"D4D5D7D9", x"DDDDD9D4", x"D3D1CECB", x"CBCAC5BF",
									 -- x"B8B4B0AF", x"AFACA8A6", x"A4A4A19F", x"A3A9ACAA", x"A5A6A8AA", x"AAA8A4A2", x"9A9B9890", x"8B8A8986",
									 -- x"8D8D8982", x"807F7C76", x"6F6B6764", x"64625C56", x"5553514F", x"4E4E4F50", x"4F535551", x"4E52585B",
									 -- x"5C595557", x"59555760", x"696F7477", x"76777B7E", x"7B818A8B", x"87827A77", x"74787B7C", x"78716F71",
									 -- x"6D6E706E", x"696B7070", x"63676567", x"6E6E6A6D", x"69696969", x"69696A6A", x"71767A7F", x"86878586",
									 -- x"848C9395", x"96979693", x"92908F90", x"92949493", x"9A9F9FA6", x"AFB5BAB3", x"B8BDC0C3", x"C3BDBCC3",
									 -- x"C7D1CEC9", x"CECCC6C8", x"D2D4D4D3", x"D4D5D3D1", x"CFD1D1CE", x"CCCDCDCD", x"D3D2D2D2", x"D1CEC9C6",
									 -- x"C4C5C5C4", x"C2C3C7CB", x"CFCED2D5", x"D3D1D0CB", x"CDC7C4C2", x"BFBFBEBA", x"B4B0AFAC", x"A7A7ACAD",
									 -- x"AEB1B2B1", x"AEADACAB", x"A5A5A5A4", x"A5A5A3A0", x"9E9C9A9A", x"98949394", x"918D8A8B", x"8B888482",
									 -- x"8E909497", x"97959290", x"908F8E8D", x"8D8C8A89", x"83838585", x"817D7C7D", x"79797A7D", x"7E7E7F81",
									 -- x"7C7A7F84", x"82828382", x"84858687", x"87868584", x"86868687", x"87888786", x"83818283", x"827E7E81",
									 -- x"7C7D7E7F", x"82848788", x"8786878A", x"8B8A8B8C", x"89888685", x"86888B8D", x"8C8B8A8C", x"91959490",
									 -- x"96969593", x"92918E8A", x"888A8987", x"8786837D", x"7C787471", x"6F6A6766", x"61616263", x"63616264",
									 -- x"61616365", x"63605F5F", x"5D5E5F5F", x"5D5A5A5B", x"5E605F5D", x"5F5E5D60", x"63646668", x"6867696B",
									 -- x"70757B7A", x"7E858894", x"A1A6ADB0", x"B0AEADAD", x"B0B5BBC1", x"C8CFD1CE", x"D0CED1D8", x"DBD9DADE",
									 -- x"E0DEDEE0", x"E2E5EAEE", x"ECEAE8E8", x"E7E7EAED", x"EFEFEEEB", x"EAEBEAE9", x"EAECECE8", x"E2DEDDDE",
									 -- x"DCDCDEE3", x"EAF0F4F5", x"F5F6F7F5", x"F4F5F7FA", x"F9F9F7F6", x"F8FAFAF8", x"F1F0F0F3", x"F4F0E7E0",
									 -- x"DBD9D7D7", x"D6D3D5DA", x"DADBDDDF", x"E0E0E1E3", x"E4E7EAEB", x"EAEAEAEA", x"E8EAEBE9", x"E6E5E8EB",
									 -- x"E8E8E9EC", x"EEF0F1F1", x"F1F2F0ED", x"EBEBE9E8", x"E9E8E7E7", x"E8E8E6E4", x"E5E4E3E4", x"E6E7E6E4",
									 -- x"E3E1DFDE", x"DFDFDFDE", x"E0E1E3E6", x"E7E8E8E8", x"E6E9EBEB", x"E9E8E9EB", x"EBE8E5E6", x"E8E8E5E2",
									 -- x"E4E2E0DE", x"DDDBDAD9", x"D6D2CFCD", x"C9C6C7CB", x"D6D7D7D7", x"DADBDAD7", x"D6D3D0CD", x"CDCBC4BE",
									 -- x"BBB5B0AD", x"ACABABAB", x"A6ABACA9", x"ACB2B1AA", x"A5A4A5A7", x"A9A8A7A7", x"9E9C9790", x"8C8B8A89",
									 -- x"8B8A8885", x"84827D78", x"746F6863", x"63615E5A", x"5753504F", x"4E4D4F51", x"4D4F5253", x"5252585D",
									 -- x"5C595556", x"59585B64", x"666F747C", x"7D7A8080", x"797B8688", x"87837B7A", x"73767472", x"7372747C",
									 -- x"7B797976", x"71727370", x"666A6D71", x"736F6B6B", x"6A6A6B6C", x"6D6F7071", x"7175787D", x"84868586",
									 -- x"86878A90", x"969A9996", x"8F929392", x"90919498", x"989B9DA9", x"B6BCBEB7", x"C1C4C2BF", x"BFBEC1CA",
									 -- x"C9CDC7C4", x"CACCC8C9", x"C8CDD2D3", x"D4D5D2CE", x"C8CACAC8", x"C8CCCDCC", x"CCCCCDCE", x"D0CFCDCA",
									 -- x"CAC7C4C5", x"C9CCCCCB", x"D2D2D5D7", x"D7D8D6CF", x"D0CDCECD", x"C9C6C3BD", x"BCB5B2B2", x"B1B4B5B2",
									 -- x"B6B8BAB9", x"B7B4B2B2", x"ACACABAA", x"A9A9A7A3", x"A3A09F9F", x"9D989697", x"98928E8E", x"8E8A8583",
									 -- x"8A8C8E8F", x"908F8D8B", x"8C8B8B8A", x"89888685", x"84828181", x"7F7B7A7A", x"7A777678", x"7A7B7C7D",
									 -- x"7A797D81", x"7F7F807E", x"80818384", x"85848483", x"83838383", x"84848382", x"817E7E80", x"807C7B7C",
									 -- x"7B7B7B7C", x"7E818385", x"84838385", x"86868789", x"87868586", x"87898A8B", x"8A8B8B8B", x"8D919291",
									 -- x"9595928E", x"8C8B8885", x"85868686", x"8684807C", x"7976726F", x"6C686564", x"63616163", x"64636160",
									 -- x"61606163", x"625F5E5F", x"5E5E5F5F", x"5D5A5B5E", x"5D605E5E", x"61616063", x"63636567", x"6767696C",
									 -- x"71747979", x"7F878A95", x"9FA3A9AE", x"B1B1B1B1", x"B0B7BFC4", x"CCD4D6D4", x"D6D5D8DD", x"DEDCDDE1",
									 -- x"E1E0E0E1", x"E3E6EBEF", x"EFF0F0EE", x"ECECECEC", x"EEEFEEEA", x"E9EAEBEA", x"E9EAEAE8", x"E2DEDCDB",
									 -- x"DCDADADE", x"E4EBF1F3", x"F4F5F6F5", x"F3F3F6F9", x"FAFAF9F8", x"F8FAFAF8", x"F2F0EFF0", x"F2F0E9E2",
									 -- x"DCDBDAD8", x"D6D6D9DB", x"DDDDE0E2", x"E2DFDFE0", x"DFE4E9EA", x"E9E8EAEB", x"EAEBEBE9", x"E8E8EAEC",
									 -- x"E9E9E9EB", x"EDF0F1F1", x"EEEFEEEB", x"EAEAE9E8", x"E9E8E7E7", x"E6E6E6E6", x"E5E4E4E4", x"E5E5E5E4",
									 -- x"E2E1E0E0", x"E0E0DFDE", x"DFE0E2E4", x"E5E6E6E6", x"E5E6E8E7", x"E6E6E7E8", x"E8E6E5E6", x"E8E9E7E5",
									 -- x"E2E1E0DF", x"DEDCDBD9", x"D5D1CFCD", x"C9C5C6CA", x"D5D5D5D4", x"D6D9D9D8", x"D4D2CFCC", x"CAC8C3BE",
									 -- x"BDB8B2AF", x"ACAAAAAB", x"A9B0B4B3", x"B2B2AFA9", x"A6A3A2A3", x"A4A3A2A4", x"9F9A9592", x"8F8C8B8A",
									 -- x"86858587", x"86817975", x"75716C67", x"64605E5C", x"59555251", x"504F4F50", x"4F4C4C51", x"5453565C",
									 -- x"5D5D5958", x"5B5B5D64", x"66727479", x"7C7D827C", x"73717B7C", x"7D7D7577", x"76766F6E", x"74777982",
									 -- x"827E7C7A", x"77787670", x"6E6E7376", x"726E6C6A", x"68696B6D", x"6F727475", x"70747577", x"7E818184",
									 -- x"8785878F", x"96969595", x"91939493", x"9192969A", x"9EA1A3AF", x"B8BCC2C1", x"C4C6C1BD", x"BEC1C4C9",
									 -- x"C8C7C5C5", x"C8CACBCA", x"C5CACECF", x"D1D4D3CF", x"CACBCBCA", x"CCD1D1CE", x"CBCBCBCD", x"CFD0CECD",
									 -- x"CCCAC8CC", x"D2D5D4D1", x"D4D5D7D6", x"D5D9D7CF", x"CECED1D2", x"CDC9C7C2", x"C2BDBCBE", x"BFC1C2BD",
									 -- x"C0C0C0C0", x"BEBBB9B9", x"B6B4B1AD", x"ABABAAA7", x"A6A3A2A3", x"A19D9C9E", x"9F989291", x"918C8786",
									 -- x"8A8A8988", x"888A8A8A", x"89888887", x"87858381", x"84807D7C", x"7B797777", x"7D797575", x"7778797A",
									 -- x"7E7B7C7E", x"7C7B7E7E", x"7B7C7E80", x"80807F7E", x"807F7F80", x"8181807E", x"827C797B", x"7C7B7A7B",
									 -- x"7C7C7B7A", x"7B7D7F81", x"82807F80", x"81828386", x"8A898888", x"88878786", x"898B8C8A", x"8A8E9192",
									 -- x"92918E8A", x"87868480", x"83828283", x"83807C7A", x"76726F6D", x"6B676565", x"67625F62", x"64635E5B",
									 -- x"605F6061", x"605E5E60", x"5F5F5F5F", x"5C5A5C60", x"5B5E5E5E", x"62636467", x"63636466", x"67696C70",
									 -- x"70727677", x"808A8E98", x"9B9EA4AA", x"AEB0B1B1", x"B0B8C1C6", x"CDD4D6D4", x"DADBDEE0", x"E0DFE0E2",
									 -- x"E1E2E3E6", x"E8E8EAED", x"EBF1F4F2", x"F1F0EEEA", x"EBEDECE8", x"E8EAEBEA", x"E9E9E9E7", x"E4DFDCDA",
									 -- x"D9D6D4D6", x"DCE4E9EC", x"F0F2F4F3", x"F1F1F4F7", x"FBFCFBFA", x"F9FAFAF9", x"F2EFEDED", x"EFEFEAE4",
									 -- x"DCDCDBD8", x"D7DADDDE", x"E0E0E3E5", x"E3DFDCDC", x"DAE0E6E8", x"E7E6E8EB", x"EDECEBEA", x"E9E9EAEB",
									 -- x"ECEBE9EA", x"ECEEEFEF", x"EAECEBE9", x"E8EAEAE8", x"EBEBEBE9", x"E7E6E8E9", x"E6E5E5E4", x"E4E4E3E3",
									 -- x"E2E1E0E0", x"E1E1E0DE", x"E0E1E2E3", x"E3E4E3E3", x"E6E5E4E4", x"E5E5E5E5", x"E6E6E5E5", x"E4E3E2E1",
									 -- x"E1E0E0DF", x"DEDDDBDA", x"D3D2D1D2", x"CEC8C6C8", x"D2D3D4D4", x"D6D8D8D7", x"D1D1CFCB", x"C8C7C4C1",
									 -- x"BCB9B6B3", x"AFA9A6A6", x"A7ADB3B5", x"B2AFAEAD", x"A6A3A2A2", x"A09D9B9B", x"9D969191", x"8F8A8787",
									 -- x"89838082", x"817C7877", x"7171706D", x"66605D5C", x"5B575454", x"53504F4F", x"5249474F", x"54525359",
									 -- x"5D5E5B59", x"5B5C5D62", x"6A777474", x"777E8479", x"77727A7B", x"7D7F787D", x"7E7B7270", x"797A787D",
									 -- x"7D79797A", x"7C7F7E76", x"74707576", x"6E6B6E6D", x"696A6A6B", x"6C6D6D6E", x"70717071", x"777A7C80",
									 -- x"84858D97", x"99959499", x"99969494", x"96989998", x"9EA0A0A8", x"ADAFBABF", x"BDC1BEBC", x"C2C6C6C5",
									 -- x"CAC8C9CC", x"CCCCCCCB", x"C9CACAC8", x"CBD2D4D1", x"CED0D0CF", x"D2D7D5D0", x"D3D1D0CF", x"CECDCAC8",
									 -- x"CACCCFD3", x"D7D9DADA", x"D6D9DBD7", x"D5D9D9D0", x"CCCCD0D0", x"CBC9C9C6", x"C4C4C9CB", x"C8C8CBC9",
									 -- x"C8C7C6C5", x"C4C1C0BF", x"BDBAB4AE", x"ACACACAA", x"ABA7A6A7", x"A6A3A2A5", x"A69D9696", x"95908C8C",
									 -- x"86868686", x"86848280", x"85848381", x"80808182", x"807F7D7B", x"79777776", x"76767575", x"75777879",
									 -- x"7B7C7A78", x"77797C7C", x"7C7B7B7D", x"7E7E7C7A", x"7A7B7C7E", x"7E7E7D7D", x"78767677", x"7879797A",
									 -- x"7D79797D", x"7D7A7B7F", x"807F7F80", x"82848484", x"81848583", x"8385888A", x"88878788", x"8B8D8B8A",
									 -- x"8C8B8986", x"8584817D", x"7A7E807F", x"7D7B7875", x"736F6C6A", x"69666667", x"66636061", x"61605F5F",
									 -- x"615E5E60", x"605F5E60", x"5F5F5F5F", x"5D5C5E61", x"5E5E6063", x"65656566", x"64686765", x"696C6D71",
									 -- x"7276797D", x"85898B8F", x"9A9B9FA6", x"ACAFB2B5", x"B4B5BAC4", x"CCCFD5DB", x"DCDBDCDF", x"E1E0E0E1",
									 -- x"E3E2E2E4", x"E7EAEBEB", x"EEF2F7F8", x"F4EFECEC", x"EAE9E7E6", x"E6E6E6E6", x"E5E7E8E6", x"E2DEDCDB",
									 -- x"D4D3D3D5", x"D6D8DDE2", x"E9EFEEE7", x"E7EBF0F5", x"FCFBFCFD", x"FBF9FAFD", x"F8F0E8E6", x"E8E9E7E4",
									 -- x"E2E0DEDC", x"DDE0E1E2", x"E4E2E2E4", x"E4E1DEDD", x"DDDFE3E5", x"E7E9EBED", x"EAE8E9EB", x"EAE7E9EE",
									 -- x"EEEBEAEA", x"EBEAECEF", x"EEEDEBE8", x"E5E6E9EB", x"ECE9E7E9", x"EAE8E7E7", x"E5E6E8E7", x"E5E2E1E0",
									 -- x"E4E1E0E1", x"E1E0E0E1", x"E0E1E1E1", x"E1E1E1E2", x"E2E3E4E5", x"E5E5E4E4", x"E2E2E2E2", x"E2E2E1E1",
									 -- x"DFDFDFDE", x"DCDAD8D6", x"D2D0D1D3", x"D4D1CDCB", x"D1D6D6D0", x"D0D6D7D1", x"CFD0CCC9", x"CAC7C3C4",
									 -- x"BEBAB5B1", x"AFADA8A3", x"AEB1B2B2", x"B3B3AFA8", x"A9A59F9C", x"9FA2A19D", x"9A96918E", x"8A858282",
									 -- x"7B7E7F7E", x"7C7C7975", x"6F6F7171", x"6D645C59", x"5C585657", x"56524D4B", x"48504B50", x"55525856",
									 -- x"5C615B54", x"595F6165", x"6275817C", x"7A7F817C", x"75777C78", x"767D7F86", x"84827E7B", x"7B7D7B77",
									 -- x"7C7D7F81", x"807B7570", x"74787A74", x"6D6A6A6B", x"6B6B6A6A", x"69696C6F", x"6E737573", x"747A7E7F",
									 -- x"8581878D", x"8D949C9B", x"94989696", x"9B99969B", x"9D9EA1A5", x"A9ACB2B6", x"BAB7BCC7", x"CDC9C7C9",
									 -- x"C8C8C8C8", x"C8C8C8C9", x"C6C8C9C8", x"C7C9CFD4", x"CDD2D6D7", x"D6D5D6D7", x"D3D4D3D1", x"D1D2D2D1",
									 -- x"C6CCCFD1", x"D5DCDFDE", x"DFDCD8D5", x"D3D2D1D0", x"CCCBCBCD", x"CDCAC9C9", x"CCCED1D4", x"D5D3D0CF",
									 -- x"CED0D1CF", x"CCCAC8C5", x"BCB7B8BA", x"B7B4B3B0", x"ACAEADAD", x"AEAAA6A8", x"AAA7A29D", x"9C99948E",
									 -- x"84838282", x"8281807F", x"81807F7E", x"7D7C7C7B", x"7A797774", x"73727273", x"73747577", x"77777675",
									 -- x"78797775", x"75787A7A", x"76787A7B", x"7B7B7B7A", x"7C7C7C7C", x"7B7A7877", x"76757473", x"74757676",
									 -- x"7876777A", x"7A777678", x"7A7A7A7D", x"80838586", x"83858583", x"82848687", x"84838286", x"8B8E8D8A",
									 -- x"8E8D8A85", x"8181807E", x"7A7D7E7C", x"79777471", x"716D6A68", x"67666668", x"65626162", x"62616162",
									 -- x"615F5E5F", x"605F5F60", x"5F5D5D5F", x"5E5D5C5D", x"5D5F6163", x"64656769", x"686C6B69", x"6E717478",
									 -- x"777B7D80", x"888B8D91", x"969AA0A4", x"A7AAADAF", x"B3B4BAC3", x"CCD1D6D9", x"D9D8D9DD", x"E0E0E1E1",
									 -- x"DFDFE0E3", x"E6E8EAEA", x"EEF1F4F4", x"F1EDEBEA", x"E5E4E2E2", x"E3E3E3E3", x"E1E1E1E0", x"E0DEDBD9",
									 -- x"D7D4D1D0", x"D0D2D7DD", x"E0E7E7E2", x"E3E9EEF4", x"FCFBFBFC", x"FBFAFAFD", x"F7F1E9E6", x"E6E7E5E3",
									 -- x"E4E5E4E1", x"E0E1E4E6", x"E5E3E3E6", x"E7E5E1DF", x"E0E1E3E6", x"E8EBEDEE", x"EBE9EAEC", x"ECEAEBF0",
									 -- x"ECEAEAEB", x"EBEAECEE", x"EDECEAE8", x"E7E7E8E9", x"EBE9E8EA", x"EBEAE8E8", x"E5E7E8E8", x"E6E4E2E1",
									 -- x"E4E2E1E2", x"E3E1E0E1", x"E0E0E0E0", x"DFDFE0E1", x"E2E3E4E4", x"E3E2E0DF", x"E2E2E2E2", x"E1E0E0E0",
									 -- x"DEDDDCDA", x"D9D8D7D7", x"D5D4D5D6", x"D4D1D0D1", x"D1D5D5D0", x"CFD3D4D0", x"CCCECBC8", x"C9C5C1C1",
									 -- x"C2C1BEB6", x"ADA6A2A1", x"A5ADB4B6", x"B4B0ACAA", x"A8A59F9A", x"999C9D9C", x"94918E8C", x"89837F7D",
									 -- x"797B7C7B", x"7A7A7875", x"71717272", x"70696462", x"57565658", x"56524F4E", x"484F4B52", x"59595D5C",
									 -- x"5E605C57", x"595D6063", x"606D7677", x"7B83837D", x"7A7B7F7A", x"787E7E83", x"82828281", x"81817D79",
									 -- x"82807D7B", x"7A787674", x"73767774", x"71707070", x"6B6A6969", x"68696D71", x"706F6E70", x"757B7D7B",
									 -- x"82808589", x"8A919998", x"97969494", x"95939397", x"9AA2A7A5", x"A4A8AFB2", x"B9B8BCC4", x"C7C5C6CA",
									 -- x"C6C7C8C9", x"C9C8C8C7", x"C7C8C9C9", x"C8CACED2", x"D5D7D9D8", x"D6D4D4D4", x"D4D2D0D1", x"D4D5D0C9",
									 -- x"CACED1D3", x"D8DEDFDC", x"E1DEDAD5", x"D2CFCCCA", x"C8C9CBCD", x"CDCDD0D3", x"D7D8DBDD", x"DDDBD8D5",
									 -- x"D5D7D7D4", x"D2CFCBC8", x"C1BBBBBE", x"BDBBBAB6", x"B3B4B1B0", x"B1ADAAAD", x"A8A6A19D", x"9B9A9590",
									 -- x"82807E7C", x"7C7D7D7D", x"7D7C7B7B", x"7C7B7877", x"76757371", x"70707071", x"70717375", x"75757473",
									 -- x"7A797673", x"74767675", x"72747677", x"76767779", x"78787979", x"78777675", x"7374726F", x"70747574",
									 -- x"71727375", x"74737170", x"77777779", x"7C7F8081", x"82848483", x"81838484", x"85828184", x"898B8885",
									 -- x"8A8B8984", x"807E7D7C", x"7A7B7B78", x"76747270", x"6F6C6968", x"67676869", x"65636263", x"63626263",
									 -- x"64626161", x"61605F5F", x"5E5C5C5F", x"615F5D5C", x"5F626565", x"6465676A", x"6A6E6E6D", x"72777A7F",
									 -- x"7D808183", x"898C8D91", x"9299A0A1", x"A2A5A8A9", x"B1B5BCC2", x"CBD4D8D9", x"D8D6D6DA", x"DDDEDEDE",
									 -- x"DADBDDDF", x"E2E5E8E9", x"ECEDEEEE", x"EDEAE9E8", x"E3E1DFDF", x"E0E1E0DE", x"DDDBD9DA", x"DDDDDAD7",
									 -- x"D5D2D0CE", x"CDCED2D6", x"D8DEDFDD", x"E0E7EEF4", x"FCFBFBFB", x"FBFAFBFC", x"F8F3ECE7", x"E5E4E3E2",
									 -- x"E4E5E6E4", x"E0DFE3E7", x"E4E2E3E6", x"E8E6E3E2", x"E3E3E4E6", x"E9ECEEEF", x"F0EEECEE", x"EDEAEAED",
									 -- x"ECEBEBEC", x"ECEBEBEC", x"EDECEBEA", x"EAE9E8E8", x"E9E7E7E9", x"EAE9E8E7", x"E6E7E9E9", x"E7E5E3E2",
									 -- x"E2E1E1E2", x"E3E1DFDF", x"E0E0E0DF", x"DEDEDFE0", x"DEDFE0E2", x"E2E1E0DF", x"E0E1E1E0", x"DEDCDCDD",
									 -- x"DCDAD8D6", x"D5D5D6D7", x"D6D7D8D7", x"D4D1D2D6", x"D1D3D2D0", x"CECECFCF", x"CACCCAC9", x"CAC7C2C2",
									 -- x"C1C0BCB5", x"ADA8A8A9", x"A9AEB6BA", x"B8B2AEAE", x"A6A4A09A", x"96969899", x"918E8A88", x"837E7A78",
									 -- x"77787978", x"77777674", x"72706F6F", x"6E6A6767", x"5B5D5F60", x"5E5A5757", x"4C504E55", x"5E606465",
									 -- x"67656360", x"5D5F6262", x"656E7577", x"7A7F7F7B", x"7B7A7D7A", x"7B808083", x"7F818382", x"82817E7B",
									 -- x"837F7A76", x"75767676", x"73747270", x"6E6E6D6B", x"6B696767", x"67686D72", x"716E6E71", x"777B7D7E",
									 -- x"80808283", x"838A9190", x"9D979697", x"93909295", x"9BA3A7A4", x"A4AAADAC", x"B2B5BABF", x"C1C0C2C4",
									 -- x"C5C6C6C7", x"C6C5C5C6", x"C7C7C8C8", x"C9CBCED0", x"D3D3D4D5", x"D4D4D4D5", x"D3D1CECE", x"D0D1CBC4",
									 -- x"C8CBCFD3", x"D9DFDFDC", x"DFDCD7D2", x"CFCCCAC9", x"D0D1D3D4", x"D2D3D7DD", x"E0E1E3E4", x"E4E2DEDC",
									 -- x"DADBDBD9", x"D7D4CFCA", x"C9C2C0C3", x"C2C2C0BB", x"BAB9B5B3", x"B4B1B0B4", x"AAA8A5A0", x"9E9C9995",
									 -- x"7F7D7B79", x"79797979", x"79777676", x"78787573", x"73727170", x"6F6E6E6E", x"6D6D6E6E", x"6F717272",
									 -- x"77757270", x"71737370", x"70717171", x"71717374", x"72727272", x"72727171", x"6D6F6F6C", x"6E737472",
									 -- x"6D6F7070", x"70706E6C", x"74747475", x"77797B7C", x"7D7F8180", x"80828383", x"84828183", x"85868481",
									 -- x"83858583", x"807E7A77", x"79797776", x"74737372", x"6F6D6A69", x"69686868", x"67666566", x"66656465",
									 -- x"67666666", x"6562605F", x"5D5C5D60", x"62615F5E", x"60636465", x"65676A6B", x"686E7070", x"75797D82",
									 -- x"83868586", x"8C8E8F93", x"91999E9D", x"9EA4A6A5", x"ADB5BCC0", x"C6D1D7D8", x"D9D5D4D6", x"D8D9D8D7",
									 -- x"D5D6D8DA", x"DCE0E5E8", x"E9E9E9E9", x"E8E7E6E5", x"E3E1DEDD", x"DDDDDBD8", x"D8D6D4D4", x"D6D6D4D1",
									 -- x"CCCDCFCF", x"CFCFD0D2", x"D3D9DADA", x"E0E7EEF5", x"FCFBFBFB", x"FBFBFAFB", x"FBF6EEE7", x"E3E2E3E4",
									 -- x"E4E5E6E4", x"E0DEE1E5", x"E2E2E2E4", x"E4E3E3E4", x"E7E5E5E6", x"E8EBEDEE", x"F2EFEDED", x"ECEAE9EA",
									 -- x"EDECECEC", x"ECECECED", x"EFEEECEC", x"ECECEBE9", x"E9E9E9EA", x"EBEAE8E7", x"E6E7E8E8", x"E8E6E4E2",
									 -- x"E1E0E0E0", x"E0DFDEDE", x"DFDFDFDE", x"DDDEE0E1", x"DCDDDEE0", x"E0E1E0E0", x"DFE0E0DF", x"DCDADADB",
									 -- x"D9D7D5D2", x"D1D2D3D4", x"D3D4D6D6", x"D3D0D1D4", x"CFCECFCE", x"CCCACCCE", x"C6C9C9C9", x"CBC8C3C2",
									 -- x"BFBAB3B0", x"B0B1B3B4", x"B7B4B3B7", x"B8B4B1B1", x"A5A3A09A", x"96939394", x"928E8883", x"7E7A7776",
									 -- x"75767575", x"74737372", x"706C6969", x"68666565", x"60616161", x"5F5C5958", x"53555458", x"60656B71",
									 -- x"726D6D6C", x"65646663", x"686F7677", x"7574777A", x"7A787A79", x"7B807E81", x"7D7F7F7D", x"7B7C7C7C",
									 -- x"7E7B7775", x"74747473", x"77777571", x"6F6F6E6D", x"6B686667", x"66666B70", x"6F6F7275", x"76777C83",
									 -- x"7F828280", x"81888D8D", x"9D95979A", x"94909495", x"9D9E9FA0", x"A6ACABA6", x"ABB0B7BC", x"BEBEBEBE",
									 -- x"C4C4C4C2", x"C1C0C2C3", x"C3C2C2C3", x"C6C9CCCD", x"CCCBCCCE", x"CFD0D2D4", x"D0CFCCC8", x"C6C7C8C7",
									 -- x"C7C9CBCF", x"D6DBDBD8", x"D9D6D1CE", x"CDCDCFD0", x"DADADBDB", x"DADADEE3", x"E4E6E7E7", x"E8E7E4E0",
									 -- x"DDDEDEDC", x"DAD8D2CD", x"CFC9C8C8", x"C5C4C3BE", x"BDBCB8B6", x"B7B5B4B8", x"B0AFABA6", x"A2A09D9A",
									 -- x"7C7A7978", x"77777575", x"75737070", x"70706F6D", x"6E6E6D6D", x"6C6A6968", x"68686869", x"6A6C6D6E",
									 -- x"6E6D6B6B", x"6D6F6F6D", x"6F6D6B6B", x"6C6E7070", x"6F6F6E6D", x"6C6B6B6A", x"696B6B6A", x"6B6F6F6D",
									 -- x"6B6C6D6C", x"6C6D6D6B", x"6E6E6F71", x"73757879", x"777A7C7D", x"7E808180", x"7D7D7F80", x"81838485",
									 -- x"8181807E", x"7F7E7974", x"77767473", x"73727273", x"6F6E6D6B", x"6A696766", x"6867686A", x"69686768",
									 -- x"67686868", x"68666360", x"605F6061", x"61605F61", x"5F606163", x"676C6D6C", x"69707475", x"7A7E8084",
									 -- x"898B8B8C", x"91929295", x"94999B9A", x"9CA3A6A4", x"A9B3BABB", x"BFCAD2D5", x"D7D3D1D2", x"D3D2D0D0",
									 -- x"D1D2D2D2", x"D4D8DEE3", x"E5E5E5E4", x"E3E2E1E0", x"E1DEDCDA", x"DAD9D7D4", x"D3D2D1CF", x"CECCCBCB",
									 -- x"C7CACDCE", x"CECECDCD", x"CFD5D7D8", x"DEE4EAF1", x"F9FAFAFA", x"FAFAFAF9", x"FBF6EFE7", x"E3E2E4E7",
									 -- x"E7E6E5E6", x"E4E1E1E3", x"E1E1E2E1", x"DFDEE1E6", x"E9E8E7E8", x"E9EBECEC", x"EDEBEAEB", x"EBEBEBEC",
									 -- x"EBEBEBEA", x"EBECEEEE", x"F0EEECEC", x"EDEDEDEC", x"EEEEEFEE", x"EEEDEBEA", x"E7E7E7E7", x"E7E5E3E2",
									 -- x"E1E0DFDE", x"DFDFDFDE", x"DDDDDDDC", x"DCDDDFE0", x"E0E0DFDF", x"DEDEDEDD", x"DEDFDFDE", x"DBD9D9D9",
									 -- x"D5D4D2D0", x"CFCFCFCF", x"CECFD1D4", x"D3D1CFCE", x"CCCBCBCB", x"CAC8C9CC", x"C3C6C5C5", x"C7C4BFBF",
									 -- x"C0BBB6B5", x"B6B6B7B9", x"BCB5B1B1", x"B1AFAFB1", x"A6A29C97", x"9391908F", x"918E8882", x"7D797674",
									 -- x"75747372", x"71706F6F", x"6C686464", x"64636364", x"66656261", x"605F5C59", x"5858595A", x"5F666E7A",
									 -- x"7B777876", x"6E6B6A64", x"64686E71", x"70707478", x"7C777977", x"797C787A", x"7C7E7E7B", x"78797A7A",
									 -- x"7B787674", x"7372706F", x"6F71716E", x"6D6E6F6F", x"69666667", x"6664676D", x"6D6E7174", x"74747A81",
									 -- x"7F838482", x"858A8F91", x"99919396", x"908E9496", x"9B97979F", x"A5A6A4A3", x"AAADB2B7", x"BABCBCBC",
									 -- x"C1C2C3C1", x"BFBDBDBE", x"BFBEBDBE", x"C1C5C7C9", x"CBC9C8CA", x"CACACCCE", x"CDCCC8C4", x"C3C5C6C6",
									 -- x"CACAC9CB", x"D0D3D3D0", x"D2D1D1D0", x"D1D3D6D7", x"DCDBDBDE", x"E0E1E4E7", x"E9EAEBEA", x"EAEBE7E3",
									 -- x"E1E2E2DF", x"DDD9D5D0", x"D2CFCFCD", x"C8C7C6C3", x"C0C0BCBA", x"BBB8B6BA", x"B4B3AFA9", x"A5A29E9B",
									 -- x"77777777", x"76757271", x"74726E6C", x"6B6B6A69", x"69696A6A", x"69676564", x"62626465", x"66676766",
									 -- x"6B6B6A69", x"696A6966", x"6A686666", x"696B6C6C", x"6D6C6B6B", x"6A6B6B6B", x"6969696A", x"6B6B6A69",
									 -- x"6A696969", x"69696A6B", x"6A6B6D6E", x"6E707172", x"73757879", x"7B7D7C7A", x"797B7C7D", x"7D7E8184",
									 -- x"84807B79", x"7A7C7974", x"75737272", x"72717171", x"70706E6C", x"6B6A6866", x"66666769", x"69676769",
									 -- x"67686969", x"6A6A6765", x"66656464", x"63616162", x"63646464", x"696E6E6A", x"6F777C7E", x"8285868A",
									 -- x"8C8F9091", x"96979698", x"999B9B9A", x"9DA3A5A4", x"A9B2B9BA", x"BDC5CED1", x"D1CFCECE", x"CECCCBCB",
									 -- x"CCCDCCCB", x"CACDD3D8", x"DDDEE0DF", x"DEDBDAD9", x"DDDCDAD9", x"D9D8D6D5", x"D0D1D1CE", x"CAC7C7C8",
									 -- x"C7CACBC9", x"C8C9CACA", x"CCD1D3D5", x"DBDFE3EA", x"F2F6F8F8", x"F8F8F9F9", x"F9F5EFE8", x"E4E4E7E9",
									 -- x"E9E6E4E6", x"E6E2E0E1", x"E1E1E1E0", x"DDDCE0E6", x"E8E9E9E9", x"E9E9EAEB", x"EAEAE9E9", x"E9E9EAEB",
									 -- x"E8E9E9E8", x"EAECEEEE", x"EEEDEBEB", x"ECEDEDEE", x"F0F1F1EF", x"EEEDECEA", x"E9E8E7E7", x"E6E5E4E2",
									 -- x"E2E2E0DF", x"DFE0E0DF", x"DBDBDBDB", x"DADBDCDE", x"DFDEDEDE", x"DDDDDDDD", x"DCDBDAD8", x"D6D5D3D2",
									 -- x"D1D0CFCE", x"CCCCCBCB", x"CCCBCCD0", x"D2D1CDCC", x"CBC9C8C8", x"C7C6C6C6", x"C3C5C4C3", x"C4C1BCBC",
									 -- x"BCBDBFBF", x"BBB6B7BB", x"B6B5B3B0", x"ABA9ACB1", x"A9A19892", x"8F8D8C8C", x"8A8A8783", x"7F7B7773",
									 -- x"74727170", x"6E6C6B6B", x"67636162", x"63636363", x"6B696562", x"6363625E", x"5A5A5C5B", x"60666E7F",
									 -- x"82838581", x"7A76726A", x"6867676B", x"6F727373", x"78737575", x"777A7678", x"797C7E7C", x"7A797876",
									 -- x"7B787471", x"706F6E6D", x"686A6A68", x"67686969", x"68656567", x"65626469", x"706E6D70", x"7376787A",
									 -- x"7F838382", x"8586878C", x"94908F8E", x"8B8D9398", x"989699A1", x"A3A0A0A5", x"A9A8A9AD", x"B0B3B7BA",
									 -- x"BBBEC1C1", x"BEBAB8B7", x"BDBCBCBD", x"C0C3C5C6", x"C7C6C6C8", x"C8C6C8CB", x"CBC8C3C2", x"C6C9C6C1",
									 -- x"C7C6C6C8", x"CBCECFCE", x"CFD1D4D7", x"D9D9DADB", x"DFDEDEE1", x"E3E5E6E8", x"ECEDEBE9", x"EAEAE7E1",
									 -- x"E2E4E3DF", x"DAD7D4D1", x"D3D2D3D1", x"CCCBCCC9", x"C5C5C2C0", x"C0BCB8BB", x"B4B3AFA9", x"A5A29D98",
									 -- x"72737374", x"7472706F", x"716F6C6A", x"68676868", x"66666767", x"67656463", x"5F606060", x"61616160",
									 -- x"66676766", x"6464625F", x"64646465", x"66676767", x"69686868", x"68696B6C", x"68656467", x"67656466",
									 -- x"68656566", x"66646568", x"68696B6B", x"6B6A6B6C", x"6E717476", x"787A7976", x"7A7A7A79", x"797A7C7F",
									 -- x"807D7875", x"76787775", x"73717073", x"74737273", x"7272706D", x"6D6E6D6B", x"69696B6C", x"6B686768",
									 -- x"6B6C6C6A", x"6B6D6C6A", x"6D6A6969", x"6A686666", x"686B6B6B", x"6E72716E", x"767E8384", x"87898B8F",
									 -- x"90959799", x"9E9E9D9E", x"A0A1A1A1", x"A1A2A4A6", x"AAB0B6B9", x"BDC3C8CA", x"CACACACB", x"CAC7C7C8",
									 -- x"C7C8C7C4", x"C0C1C5C9", x"D1D5D9DA", x"D9D6D5D4", x"D6D7D7D6", x"D5D4D3D4", x"CCCDCECC", x"C8C6C6C6",
									 -- x"C6C8C9C6", x"C5C7C9C9", x"CBD0D2D5", x"DADCDFE5", x"EAF0F5F5", x"F5F6F8F8", x"F8F5F0EB", x"E9E9EAEC",
									 -- x"E8E4E3E6", x"E5E1DEDE", x"DFDEDDDE", x"DDDDDFE2", x"E2E5E8E8", x"E7E5E6E8", x"EBEBEBEA", x"E8E8E9EA",
									 -- x"E9EBEBEA", x"EAECEDEC", x"EBECECEC", x"ECEDEEF0", x"EFF1F0EE", x"ECECEBE9", x"ECEBE9E8", x"E7E7E5E4",
									 -- x"E1E2E1DF", x"E0E1E1DE", x"DCDCDCDC", x"DBDBDBDC", x"DADBDCDD", x"DDDCDBDB", x"DAD8D5D3", x"D2D0CCCA",
									 -- x"CCCCCBCA", x"C9C9C8C8", x"CAC8C8CB", x"CECECDCD", x"CCCAC7C4", x"C4C4C2BF", x"C3C4C2C0", x"C2BFBBBC",
									 -- x"BABBBFC1", x"BDB7B8BD", x"B5B6B4AE", x"A9A8ABAE", x"A9A29994", x"908B8988", x"86878581", x"7E7B7671",
									 -- x"72706E6E", x"6C696868", x"66636265", x"68676665", x"69696562", x"6162615F", x"5E5C6161", x"656A6D7D",
									 -- x"858E8F89", x"86827A72", x"6E6C6A6A", x"6D70706E", x"716C7071", x"74767376", x"75797C7C", x"7A797572",
									 -- x"7673706D", x"6D6C6C6B", x"6C6C6B69", x"696A6866", x"68646366", x"64606267", x"6D6E6D6D", x"6F737575",
									 -- x"7A7E7D7F", x"827E7D85", x"8E918F8B", x"8B8D9094", x"9596999E", x"A09FA0A3", x"A5A1A1A5", x"A6A7ADB5",
									 -- x"B5B9BBBB", x"B8B5B4B4", x"B7B8BABC", x"BFC1C3C4", x"C1C0C2C5", x"C4C2C3C8", x"C7C4C1C1", x"C5C7C3BD",
									 -- x"C0C0C2C5", x"C8CBCDCE", x"CED1D5D9", x"DBDCDEDF", x"E6E5E5E6", x"E5E4E6E9", x"EAEBEAE7", x"E8E9E6E0",
									 -- x"E0E2E2DD", x"D8D5D5D4", x"D3D2D4D2", x"CFCFCFCB", x"C8C8C5C4", x"C4BFBCBE", x"B8B5B0AB", x"A7A29B95",
									 -- x"6F6F7071", x"72716F6E", x"6A6A6967", x"65656566", x"63636364", x"63636262", x"615F5D5B", x"5B5C5E5F",
									 -- x"595D5F5F", x"5F5F5E5D", x"61636565", x"64626263", x"67666463", x"62626364", x"625D5C61", x"615E5E63",
									 -- x"67626265", x"65616164", x"62646769", x"696A6B6C", x"6A6D7174", x"76787775", x"79787676", x"77797B7D",
									 -- x"78787674", x"74757574", x"71707074", x"76767676", x"7575726F", x"6F727371", x"71717272", x"706C6A6B",
									 -- x"71716F6C", x"6C6E6F6E", x"726E6C6E", x"71706D6B", x"686D7071", x"73797A78", x"7A828586", x"898B8D91",
									 -- x"979C9FA2", x"A8A7A5A6", x"A5A6A8A8", x"A5A3A5A9", x"A8ABB0B5", x"BBBFC1C2", x"C7C7C9CA", x"C7C4C4C6",
									 -- x"C3C5C4C0", x"BBB9BBBF", x"C7CDD3D7", x"D6D4D3D3", x"CFD0D2D0", x"CECDCDCE", x"C6C7C8C7", x"C5C3C3C3",
									 -- x"C3C6C7C6", x"C6C9CBCB", x"CDD1D4D6", x"DBDDDFE4", x"E4EBF2F3", x"F3F5F7F8", x"F8F5F2EF", x"EEEEEEEF",
									 -- x"E8E5E5E7", x"E6E0DEDF", x"DEDBDADC", x"DEDEDEDE", x"DDE1E5E6", x"E3E2E3E5", x"E8EAEBEA", x"E9E9EBED",
									 -- x"EDEFEFED", x"ECEDEBE9", x"EBECEDEE", x"EDEEF0F1", x"F0F2F1EE", x"ECEDECEA", x"EFEDEAE9", x"E8E8E7E6",
									 -- x"DFE1E1DF", x"E0E1DFDD", x"DEDFDFDE", x"DCDCDCDC", x"DADBDCDD", x"DCD9D6D5", x"DCD8D5D3", x"D2CFCBC7",
									 -- x"C9C9C8C8", x"C7C7C7C6", x"C9C6C5C7", x"C9CBCDCF", x"CDCCC7C3", x"C2C3BFBA", x"BFC0BDBC", x"BEBDBABC",
									 -- x"BDBAB9BB", x"BBB8B8BA", x"B8B6AFA8", x"A7AAAAA8", x"A7A29D99", x"938C8684", x"8786837E", x"7A787470",
									 -- x"706E6C6C", x"6A676667", x"6B69696C", x"6E6D6B69", x"6E6F6D68", x"65656564", x"63606666", x"6A6E6C7A",
									 -- x"8391928B", x"8A887C74", x"6C6E6D69", x"67696C6D", x"6F6B6E6E", x"70716D70", x"73767777", x"77767370",
									 -- x"6F6D6B6B", x"6B6B6A69", x"69686666", x"696A6763", x"67636264", x"635F6167", x"666C6E6A", x"686B7073",
									 -- x"7276777C", x"827C7B86", x"8791908B", x"8C8C8A8C", x"92929397", x"9DA1A09C", x"A19E9FA4", x"A3A0A6B1",
									 -- x"B3B4B5B3", x"B0AFB1B3", x"ACAFB4B8", x"BBBDBFC0", x"BDBDC0C2", x"C0BBBCC1", x"C2C2C2C0", x"C0C1C0BF",
									 -- x"BDBEC0C3", x"C6C7C9CA", x"CDCFD2D5", x"D8DCE1E4", x"E6E6E7E7", x"E4E4E7EC", x"E9EBE9E7", x"E8EAE7E1",
									 -- x"E0E2E2DE", x"D9D8D9DB", x"D3D2D3D2", x"D0D1D0C9", x"C7C8C5C4", x"C5C1BFC1", x"BDBAB3AD", x"A9A39B93",
									 -- x"74727070", x"706F6B68", x"67666462", x"60606263", x"605F5E5D", x"5D5D5D5D", x"5C5A5859", x"5B5B5957",
									 -- x"5956575C", x"5D59585A", x"5D5E5E5F", x"6162615F", x"62626161", x"61606060", x"5C5D5E5F", x"5F5E5D5C",
									 -- x"5E5E5E5E", x"5F606263", x"5E5F6163", x"65686A6B", x"6B6A6C71", x"74737170", x"73717173", x"76777879",
									 -- x"77797874", x"7171716F", x"74747574", x"72727476", x"77767474", x"76767573", x"7A777372", x"73737270",
									 -- x"70736E70", x"696F6E71", x"6F716F6D", x"71727274", x"71707075", x"7A77777E", x"8183878C", x"8F909499",
									 -- x"9EA0A0A5", x"ABABABAF", x"ABABAAA9", x"A8A8A9AA", x"ADAEAFAF", x"B1B7BCBF", x"C1C2C5C8", x"C5C0C0C3",
									 -- x"C2BDBDBF", x"BAB3B6BF", x"BDC2C7CB", x"CCCCCCCC", x"C9CACBCA", x"CAC9C9CA", x"C5C7C6C3", x"BFBEBFC1",
									 -- x"C0C1C4C6", x"C7C8C8C8", x"CACED1D3", x"D5DADDDE", x"E0E2E8EF", x"F3F3F3F5", x"F5F6F5F2", x"F0F0F0F0",
									 -- x"EBE8E4E0", x"DEDCDAD8", x"D9DADBDB", x"DAD8D7D7", x"DADEE3E5", x"E4E1E0DF", x"E9E8E6E6", x"E8EAEBEC",
									 -- x"F0F1F0EE", x"EEF0EFEC", x"EFEFEFEF", x"EEEEEDED", x"F0F2F2F0", x"EDEBECED", x"ECECEAE6", x"E5E6E7E6",
									 -- x"E3E2E1E1", x"E0DFDDDC", x"DDDCDCDD", x"DEDDDCDA", x"DBD9D8D9", x"DAD8D7D7", x"D6D3D0CE", x"CDCBC7C4",
									 -- x"C8C8CACC", x"CAC7C5C6", x"C7C5C6C9", x"CAC9CACD", x"CBCAC7C5", x"C4C2BEB9", x"BEBBBABC", x"BCB9BABD",
									 -- x"B7B8B9BA", x"B9B9B8B7", x"B4B4B0AB", x"A8A6A4A2", x"A3A09E9C", x"99928A84", x"85817C7A", x"7A797774",
									 -- x"70736C6A", x"706C676F", x"6A737272", x"77716A72", x"6D70726C", x"63636766", x"6469696E", x"7571727E",
									 -- x"80888E8D", x"86817E7C", x"726D6D6F", x"6C6B6C6B", x"67696C6F", x"706F6E6D", x"6E717374", x"74727171",
									 -- x"6C706B68", x"696B6C64", x"68666361", x"63666663", x"63626465", x"6562605F", x"62666969", x"67676B6E",
									 -- x"7374777C", x"7D7C7D7F", x"82868A8D", x"908F8B85", x"8A8A8E95", x"9A9A9A9D", x"9D9FA09D", x"9C9FA6AB",
									 -- x"ADADAEAE", x"ACAAABAD", x"A9B2B3AE", x"B1B8BABA", x"BCBBB9B7", x"B7B9BCBE", x"C0BFBDBB", x"BDBFBFBD",
									 -- x"BBB5B8C3", x"C5BFC1CC", x"D0D0D4DA", x"DDDFE2E5", x"E8E6E5E5", x"E5E4E6E8", x"E6E8E8E5", x"E3E4E4E4",
									 -- x"E4E0DDDE", x"DDD9D6D6", x"D5D8D9D6", x"D3D1CFCD", x"CBCBC8C4", x"C4C5C3C0", x"C2BCB4AD", x"A8A19890",
									 -- x"706E6D6C", x"6C6B6967", x"66656361", x"5F5E5D5D", x"5B5B5B5A", x"5A5A5A5A", x"59575656", x"57575553",
									 -- x"5A565659", x"59575759", x"5B5B5A59", x"595A5957", x"5D5D5C5C", x"5C5C5B5B", x"5657585A", x"5B5B5B5A",
									 -- x"5B5B5B5B", x"5B5C5D5D", x"5D5D5F60", x"62656667", x"6766676B", x"6E6E6E6E", x"716F7073", x"75757576",
									 -- x"7A747274", x"716C6F75", x"77767575", x"76777878", x"7A797879", x"7A7A7978", x"78777676", x"76777877",
									 -- x"77787374", x"6F737275", x"7677726D", x"6F717275", x"79787678", x"7B7B7C82", x"84868B8F", x"9092989E",
									 -- x"9EA1A3A7", x"ACADAFB4", x"B4B3B2B0", x"AEADADAD", x"AEB0B0B0", x"B2B7BCBE", x"BDBFC3C6", x"C5C2C0C0",
									 -- x"BFB9B6B7", x"B4AFAFB3", x"B7BABEC0", x"C0BFBFC0", x"C5C6C7C5", x"C3C2C3C4", x"C2C3C2BF", x"BCBDC0C3",
									 -- x"C1C1C1C3", x"C5C7C7C7", x"C8CCCFD0", x"D3D9DEE0", x"E2E3E7EC", x"F0F0F1F3", x"F6F6F4F2", x"F2F4F5F5",
									 -- x"EDEAE5E1", x"DDD9D5D3", x"D5D6D6D6", x"D5D5D5D5", x"D9DCDFE3", x"E4E3E1E0", x"E3E3E4E5", x"E7EAECED",
									 -- x"EEEFEFED", x"EEF0EFED", x"EFF0F0EF", x"EFEFEFEE", x"EFF0F0EF", x"ECEBEBEC", x"ECEBE9E6", x"E5E5E5E4",
									 -- x"E3E2E1E0", x"DFDEDCDB", x"DCDBDADA", x"DADAD9D9", x"D8D6D5D7", x"D8D7D5D5", x"D5D2CFCC", x"CAC8C6C4",
									 -- x"C8C8CACB", x"CAC8C7C8", x"C6C4C3C5", x"C6C6C7CA", x"C9CAC9C6", x"C3C0BCB8", x"BAB8B8BA", x"B8B5B6BA",
									 -- x"B7B8B8B7", x"B7B7B7B7", x"B4B4B0AB", x"A8A6A5A2", x"9F9E9D9E", x"9C97908A", x"85837F7B", x"78757372",
									 -- x"6F727172", x"76726F74", x"777E7976", x"7B766F74", x"7473736F", x"67666865", x"666B6E74", x"7D7E7F88",
									 -- x"82878B87", x"7D78797D", x"756F6E6E", x"6A696A69", x"686A6C6E", x"6F6E6D6C", x"6B6D7070", x"6F6D6C6D",
									 -- x"6A6E6B6C", x"6A65645F", x"63615F5E", x"6063625F", x"5F5D5B5C", x"5C5C5E60", x"62656869", x"68686A6C",
									 -- x"6C6D7175", x"78787B7E", x"8385878B", x"8F908C86", x"86878C92", x"96979797", x"9C9D9E9D", x"9B9CA1A5",
									 -- x"A5A6A9AA", x"A9A7A7A9", x"ABADACAE", x"B3B6B6B8", x"B6B6B4B3", x"B3B5B8BA", x"BBBBB9B8", x"BABCBCBA",
									 -- x"B7B7BBC1", x"C4C2C5CA", x"D1D2D6DB", x"DDDEDFE2", x"E5E3E3E4", x"E4E3E4E6", x"E4E4E4E3", x"E4E4E2DF",
									 -- x"E2DEDCDC", x"DBD7D4D2", x"D4D5D4D2", x"D1D0CECB", x"CCCBC9C6", x"C5C6C4C1", x"BEB8B1AC", x"A8A29B95",
									 -- x"6D6D6C6C", x"6B6A6868", x"65646462", x"605E5C5B", x"58585757", x"57565656", x"54545353", x"53535252",
									 -- x"59555354", x"54535558", x"57575655", x"55575756", x"58585858", x"59595958", x"54555758", x"595A5A5A",
									 -- x"59595959", x"59595A5A", x"5A5B5C5D", x"5F606162", x"64646467", x"696A6C6F", x"6E6D6E72", x"73737273",
									 -- x"75706F72", x"716E7077", x"79777676", x"797A7A7A", x"7A7B7C7C", x"7D7C7C7B", x"78787979", x"797A7B7C",
									 -- x"7B7A7677", x"74767576", x"797B7771", x"71727477", x"787A797A", x"7F818387", x"85888E91", x"919399A0",
									 -- x"9FA3A6A9", x"AEB1B5BC", x"BFBEBCBA", x"B7B5B3B1", x"B4B5B5B4", x"B5B8BBBC", x"BABDC1C4", x"C7C7C3BE",
									 -- x"BFB9B4B3", x"B3B1ADAA", x"B3B5B7B8", x"B7B7B7B8", x"BCBEBEBC", x"B9B8BABC", x"C0BFBDB9", x"B6B6B9BD",
									 -- x"C0C0BFC0", x"C2C5C6C7", x"C8CACDCE", x"D2D7DDE0", x"E3E3E6EA", x"ECEDEFF2", x"F4F5F4F4", x"F6F8F7F5",
									 -- x"EFECE8E4", x"DFD9D4D0", x"D1D0D0D1", x"D2D3D5D6", x"D6D7DADE", x"E2E3E2DF", x"DDE0E3E5", x"E7E9EBED",
									 -- x"EDEDEDED", x"EEF0F0EE", x"EFEFEFEF", x"EFEFEFEF", x"EEEEEEEE", x"EDECECEB", x"EBECEAE6", x"E5E5E5E3",
									 -- x"E3E1E0DF", x"DDDCDAD9", x"D9D9D8D7", x"D6D6D6D7", x"D5D3D2D4", x"D5D4D3D3", x"D2CFCBC7", x"C4C3C3C3",
									 -- x"C6C6C8CA", x"C9C7C7C8", x"C6C4C3C3", x"C3C4C6C8", x"C5C8C8C4", x"C0BCB9B6", x"B8B7B8B9", x"B8B5B5B8",
									 -- x"B7B6B5B5", x"B4B4B4B5", x"B2B1AFAA", x"A7A6A4A2", x"9B9A9B9C", x"9B98918B", x"8584817C", x"76727070",
									 -- x"6D71767A", x"7C7C7D80", x"898D847C", x"7F7D7676", x"7A747270", x"6B696968", x"686D7179", x"8488888B",
									 -- x"86817D7D", x"7D797778", x"736D6B6A", x"67666766", x"67696B6C", x"6C6B6A69", x"686B6E6E", x"6C6A6A6C",
									 -- x"70727072", x"6D636261", x"5E5D5B5A", x"5C5E5C5A", x"59595A5D", x"5E5D5D5E", x"60626567", x"6868696A",
									 -- x"68696C70", x"7275787C", x"7F808286", x"8C8F8C87", x"84888C90", x"93959594", x"9998999A", x"99989A9E",
									 -- x"A0A0A2A4", x"A4A3A5A8", x"ABA5A1A7", x"AFAFAEB4", x"B1B1B0B0", x"B0B1B3B5", x"B5B5B4B4", x"B6B8B8B6",
									 -- x"B6BCC1C3", x"C6CBCCCB", x"D0D2D6DA", x"DCDCDDDE", x"E0DFE0E2", x"E3E2E1E2", x"E1E0DFE0", x"E2E3DFD9",
									 -- x"DEDCDADA", x"D9D6D4D2", x"D6D5D3D1", x"D1D2D0CC", x"CCCBC9C7", x"C7C7C5C2", x"BCB6AFA9", x"A5A09994",
									 -- x"696A6C6C", x"6A686767", x"62616160", x"5F5E5D5B", x"59585655", x"53535353", x"50505151", x"51525252",
									 -- x"55524F50", x"50505254", x"53545453", x"54565755", x"53535354", x"56575757", x"56565757", x"58585858",
									 -- x"58585858", x"59595958", x"58595A5B", x"5C5D5E5E", x"62626265", x"66676A6D", x"6C6C6D70", x"71717071",
									 -- x"6C707271", x"71747574", x"79787777", x"787A7A7A", x"7D7E8081", x"807F7F7F", x"7B7B7A79", x"79797979",
									 -- x"7C7A7779", x"79797778", x"767B7B79", x"79797779", x"777C7D7E", x"83868586", x"888B8F91", x"93969CA1",
									 -- x"A1A6A8AB", x"B2B6BBC2", x"C6C5C4C2", x"C0BDBAB8", x"BBBCBCBA", x"BABCBDBC", x"BDBFC2C5", x"CACDC8C0",
									 -- x"C1BDB7B5", x"B5B4AFA9", x"B0B1B3B4", x"B5B5B7B7", x"B5B7B8B6", x"B4B3B5B8", x"BAB9B8B6", x"B4B2B4B7",
									 -- x"BCBDBFC0", x"C0C2C5C7", x"C8CACDCF", x"D2D6DBDE", x"E1E2E5E8", x"EAECEFF2", x"F2F3F6F7", x"F9F9F5F0",
									 -- x"EFEDEAE7", x"E3DDD7D2", x"CFCFCFD0", x"D2D4D6D7", x"D3D4D6DA", x"DEE0E0DE", x"DBDEE3E5", x"E6E7E9EB",
									 -- x"ECEDEDEE", x"EFF1F1F0", x"EEEEEEEE", x"EEEEEFEF", x"EFEFEFEF", x"EFEFEEED", x"ECECEBE8", x"E6E6E4E3",
									 -- x"E2E1DFDD", x"DCDAD9D7", x"D6D7D7D7", x"D5D4D5D6", x"D5D3D1D3", x"D3D1D0CF", x"CDCBC7C3", x"BFBDBEBF",
									 -- x"C2C3C5C8", x"C8C6C5C6", x"C5C4C3C2", x"C1C2C3C4", x"C2C3C3BF", x"BCBAB6B3", x"B7B6B6B8", x"B9B7B6B7",
									 -- x"B4B4B3B2", x"B2B1B1B1", x"ADAEACA8", x"A6A5A4A2", x"9D9C9A9A", x"99968F89", x"8684807B", x"7672706F",
									 -- x"6E727C83", x"85898F92", x"96978D81", x"80807B79", x"79716E6F", x"6C6B6E6F", x"676B7179", x"858C8C8A",
									 -- x"897F797C", x"7E797371", x"6D696868", x"65656664", x"64656768", x"68676665", x"64676B6C", x"6A696A6C",
									 -- x"70716C6B", x"665F605F", x"5E5C5B5A", x"5A5A5856", x"5A5A5D60", x"615F5E5E", x"5E5F6063", x"66686968",
									 -- x"66676A6C", x"6D707477", x"77797C81", x"868B8A88", x"84898C8D", x"90949593", x"96939497", x"98959497",
									 -- x"9C9B9A9B", x"9C9DA1A5", x"A8A19A9F", x"A7A8AAB1", x"AEAFAFAE", x"ADAEAFB0", x"AFB0B1B1", x"B3B5B5B4",
									 -- x"B7BEC4C7", x"CACFD0CE", x"CFD0D4D7", x"D9DADBDC", x"DDDDDFE1", x"E2DFDEDE", x"DFDEDDDC", x"DEDFDBD5",
									 -- x"D9D7D5D5", x"D5D4D3D3", x"D7D6D3D0", x"D0D1D0CE", x"CBCAC8C7", x"C7C6C3C1", x"B8B2ABA6", x"A29C9692",
									 -- x"6366696A", x"68666464", x"5F5E5C5B", x"5B5A5959", x"5A585552", x"504F4F4F", x"4D4E4E4F", x"4F505051",
									 -- x"4F4D4C4C", x"4D4E4F50", x"4F515251", x"5051504F", x"504F4F50", x"52545352", x"54545453", x"53535454",
									 -- x"55545456", x"57585757", x"5657585A", x"5B5C5C5D", x"5E5E5F62", x"63636567", x"6B6B6C6E", x"6F6F7071",
									 -- x"6C707372", x"72747573", x"76777878", x"797A7D7F", x"84858788", x"87878686", x"827F7C7B", x"7B7C7A78",
									 -- x"7D7A7B7D", x"7F7D7C7C", x"787E7F7F", x"81807E7F", x"7F838383", x"86878586", x"8D8F9194", x"979CA1A3",
									 -- x"A5A8A9AC", x"B5BBBFC4", x"C7C7C6C6", x"C6C4C1BF", x"C0C1C1C0", x"C0C1C1C0", x"C3C4C4C6", x"CBCFCBC4",
									 -- x"C0BEBAB6", x"B5B5B1AC", x"AEAFB1B3", x"B4B4B5B6", x"B4B5B6B5", x"B2B2B4B7", x"B2B2B3B5", x"B5B3B4B6",
									 -- x"B6BBBFC0", x"BFBFC3C7", x"C7C9CDD0", x"D3D6D9DC", x"DCDFE4E7", x"EAEDF0F2", x"F2F3F5F7", x"F9F8F3EE",
									 -- x"EEEDEBE9", x"E6E0DAD6", x"D3D2D1D1", x"D3D4D4D4", x"D1D3D6D8", x"DBDCDCDD", x"D9DDE1E4", x"E5E5E7E9",
									 -- x"EBEBECEF", x"F0F1F1F1", x"EFEEEEEE", x"EEEEEEEE", x"EFEFEFF0", x"F0F0EFEE", x"EAEBEBE8", x"E6E6E4E1",
									 -- x"E2E0DEDC", x"DAD9D7D6", x"D4D6D7D8", x"D6D5D4D5", x"D6D3D2D2", x"D1CFCDCC", x"CAC8C5C1", x"BDBBBBBC",
									 -- x"BFC0C4C8", x"C8C5C4C4", x"C1C1C0BF", x"BEBEBEBD", x"C0BFBDBA", x"BAB9B6B3", x"B4B2B2B5", x"B7B7B4B2",
									 -- x"B1B1B1B1", x"B0AEADAC", x"AAAAA9A7", x"A5A5A5A3", x"A2A09C9A", x"9998928C", x"88847F7A", x"7673716F",
									 -- x"7077848D", x"8F949A9B", x"9A9A9185", x"80807F7C", x"77706F70", x"6F707678", x"6C6D737C", x"878F908B",
									 -- x"8682807F", x"776D6B6F", x"6A686868", x"66666763", x"61626364", x"65646463", x"61646767", x"66656668",
									 -- x"6C6F6964", x"6160625C", x"5E5C5B5B", x"5B595756", x"5D5A595A", x"5B5C5E61", x"605F5E60", x"64676767",
									 -- x"63656868", x"686B6E71", x"71757A7D", x"80848685", x"83878A89", x"8B909392", x"94939396", x"96939293",
									 -- x"96959596", x"97989B9E", x"A1A09C9D", x"A3A6A8AC", x"A9AAAAAA", x"AAAAAAAB", x"ACAEAFAF", x"B1B4B4B3",
									 -- x"B6BAC0C5", x"C8CACBCC", x"CFD1D2D4", x"D5D7D9DA", x"DADADCDF", x"DFDCDADA", x"DCDCDBD9", x"D8D8D6D4",
									 -- x"D3D2D0CF", x"CFD0D1D1", x"D1D2D1CE", x"CCCDCFCF", x"CBCAC8C7", x"C6C4C1BF", x"B3ADA7A4", x"A09B9694",
									 -- x"60636668", x"66646261", x"605D5A58", x"58575655", x"5755524F", x"4C4B4B4C", x"4C4B4B4B", x"4C4C4B4B",
									 -- x"4A494949", x"4A4B4B4B", x"494C4D4D", x"4D4E4E4C", x"504F4D4E", x"5151504F", x"51505050", x"50515252",
									 -- x"53525254", x"56575757", x"54555758", x"5A5B5B5B", x"5C5C5D61", x"62626263", x"68686A6C", x"6D6D6E70",
									 -- x"736F7074", x"736F7178", x"76787A7B", x"7C7E8285", x"88898A8C", x"8C8C8C8C", x"89868181", x"8283817F",
									 -- x"817D8081", x"85808181", x"81858584", x"87888687", x"86878584", x"8788888C", x"8F919395", x"9AA0A3A4",
									 -- x"A8ABAAAD", x"B6BDC0C4", x"C6C6C7C9", x"CACAC8C6", x"C3C5C6C6", x"C8CAC9C7", x"C8C8C6C7", x"CBCDCAC6",
									 -- x"C0C0BEBA", x"B8B6B4B2", x"B0B0B1B2", x"B3B3B3B3", x"B2B3B3B2", x"B0B0B1B2", x"B0AFB0B3", x"B3B0B0B2",
									 -- x"B3B8BEBF", x"BDBDC0C4", x"C3C6CBD0", x"D3D5D8DA", x"D7DCE2E5", x"E8ECEFF1", x"F2F3F3F3", x"F4F5F3F0",
									 -- x"ECEBEAE8", x"E6E1DCD8", x"D7D5D2D1", x"D1D1D0CF", x"D2D3D5D6", x"D7D8D9D9", x"D5D8DCDF", x"E1E2E4E6",
									 -- x"E8E8EAEE", x"F1F1F1F1", x"F0EFEFEE", x"EEEEEEEF", x"EDEDEEEF", x"EFEEEEED", x"E9EAEAE8", x"E7E6E3E1",
									 -- x"E1E0DDDB", x"D9D8D7D6", x"D4D5D7D8", x"D7D5D3D3", x"D6D3D1D1", x"D0CDCBCA", x"C8C6C3C0", x"BEBCBCBC",
									 -- x"BEBFC3C6", x"C7C4C2C2", x"BFBFBFBD", x"BCBCBBBA", x"BEBCB9B7", x"B8B9B6B3", x"B2B1B2B4", x"B7B6B3B0",
									 -- x"AEAFAFAE", x"ADABA9A8", x"A8A9A8A6", x"A5A6A5A4", x"A09E9A97", x"999A968F", x"8A86807B", x"77757371",
									 -- x"737E8A92", x"96989899", x"9A989289", x"83828280", x"7A747375", x"757A7F81", x"7D787B82", x"888D8D86",
									 -- x"817D7A77", x"716B6A6D", x"68666766", x"6364645F", x"60616162", x"62626262", x"61636464", x"63636363",
									 -- x"666C6864", x"6363645B", x"5C5B5A5B", x"5B595858", x"57565658", x"595A5C5E", x"62605E5F", x"61646464",
									 -- x"61656867", x"67696C6F", x"6E73787A", x"7B7D8081", x"84868787", x"888C8F91", x"93939495", x"94939190",
									 -- x"92929395", x"97969798", x"959B9C9C", x"A0A3A3A3", x"A1A2A4A4", x"A5A6A7A8", x"ABADAEAE", x"AFB2B3B3",
									 -- x"B5B7BCC2", x"C5C4C5C9", x"CFD1D1D1", x"D1D3D5D5", x"D6D6D8DB", x"DAD8D6D6", x"D7D9D8D4", x"D2D2D2D2",
									 -- x"D2D2CFCD", x"CCCDCECE", x"CCCFCFCD", x"CCCDD0D1", x"CBC9C7C7", x"C5C1BDBB", x"B2ACA6A3", x"9E979290",
									 -- x"5F616363", x"6361605F", x"605D5A57", x"57565452", x"51504E4D", x"4B4A4A49", x"49484747", x"49494847",
									 -- x"47474747", x"48484847", x"44474949", x"494B4C4C", x"4F4D4C4D", x"5051504E", x"4F4F4E4E", x"4F505152",
									 -- x"51504F51", x"54565655", x"52535557", x"58585958", x"5A595A5E", x"61616161", x"6364676A", x"6B6A6B6D",
									 -- x"716D6F74", x"74707278", x"797A7B7D", x"7F828587", x"8A898A8C", x"8E90908F", x"918E8A89", x"8A8B8C8B",
									 -- x"8A858886", x"89838788", x"8B8D8B8A", x"8F908E8E", x"8A898788", x"8C8C8D93", x"8F929597", x"9BA1A4A5",
									 -- x"A9ADADAE", x"B5BBBFC3", x"C7C7C8CB", x"CECFCDCB", x"C9CBCDCE", x"D1D2D1CE", x"CDCBC9CA", x"CAC8C7C7",
									 -- x"C4C3C1C0", x"BDBAB9BA", x"B5B4B2B2", x"B2B2B2B2", x"AFAFAFAF", x"AFAFAFAF", x"B4B1B0B1", x"B0ADADB0",
									 -- x"B3B6BABC", x"BCBCBDBF", x"C1C3C8CE", x"D1D1D4D7", x"D4DADFE1", x"E4E8ECEE", x"F0F0F0EE", x"EEEFEFEE",
									 -- x"E9E8E7E7", x"E6E3DFDC", x"D9D6D2D0", x"CFCFCECD", x"D2D1D0D1", x"D3D4D4D3", x"D2D3D5D8", x"DBDDDFE0",
									 -- x"E2E2E6EC", x"F0F0F0F0", x"F0F0EEED", x"EDEDEDED", x"EBEDEFEF", x"EEECECED", x"E9EBECEA", x"E9E8E5E2",
									 -- x"E1DFDCDA", x"D9D8D7D6", x"D5D5D5D6", x"D5D4D2D0", x"D2D0CECF", x"CECCCAC9", x"C5C3BFBD", x"BDBDBDBC",
									 -- x"BDBEC0C3", x"C2C0BFC0", x"BEBEBDBA", x"B9BAB9B8", x"B9B9B7B6", x"B5B6B4B1", x"B1B3B6B7", x"B7B5B2B0",
									 -- x"AEADADAC", x"AAA8A7A6", x"A5A7A6A4", x"A3A4A3A1", x"9C9A9794", x"9699948D", x"8986817C", x"77767677",
									 -- x"7C899094", x"9A9A979A", x"9A95918D", x"88878683", x"7E79797B", x"7E868986", x"887E7D83", x"8384847E",
									 -- x"7B77726F", x"6D6C6A68", x"65646462", x"5F61615C", x"60606060", x"5F5F5F5F", x"5F5F6060", x"60605F5E",
									 -- x"5D636261", x"5F5B5C57", x"5A585859", x"58575657", x"53545659", x"5A595858", x"5E5C5B5C", x"5E606160",
									 -- x"60656868", x"67686A6B", x"6B6F7273", x"74787B7C", x"84848586", x"8686898D", x"8D919290", x"8F91918F",
									 -- x"908E8E90", x"92929395", x"8F959798", x"9D9F9C9C", x"9FA0A1A2", x"A3A4A6A7", x"AAACACAC", x"ADB0B2B2",
									 -- x"B6B7BABF", x"C0C0C2C5", x"CACCCDCC", x"CDCFD0D0", x"D1D1D3D5", x"D5D3D2D2", x"D1D3D2CF", x"CDCDCECE",
									 -- x"CECFCECB", x"CACBCCCB", x"CBCDCDCC", x"CCCECECE", x"CAC7C5C4", x"C2BCB7B5", x"B2ABA5A1", x"9B928B8A",
									 -- x"5D5D5D5E", x"5E5D5C5B", x"5D5A5755", x"5554514F", x"4C4D4D4D", x"4C4B4A49", x"47454445", x"48494846",
									 -- x"46464645", x"46464645", x"45474745", x"44454646", x"4A484749", x"4D4F4E4D", x"4E4E4D4C", x"4C4D4E4F",
									 -- x"4E4C4B4C", x"4F515251", x"51525455", x"56575656", x"5655565A", x"5E5F5E5E", x"5F616569", x"6968696A",
									 -- x"686D7172", x"73767675", x"7D7C7C7D", x"81848585", x"8A8A8A8C", x"90939392", x"9593918F", x"8F909294",
									 -- x"948E908C", x"8F878D90", x"8F919090", x"96979392", x"918F8E91", x"94908F95", x"90969A9C", x"9EA3A7A9",
									 -- x"A8AEB0AF", x"B4B9BDC3", x"C8C8C9CD", x"D0D1D0CE", x"D0D2D4D5", x"D7D8D6D3", x"D0CDCCCD", x"CAC6C5C8",
									 -- x"C7C4C3C2", x"C0BCBBBD", x"B7B5B2B0", x"B0B0B1B2", x"AFAEAEB0", x"B2B3B2B1", x"B8B3B1B2", x"B2B1B3B8",
									 -- x"B4B5B7B9", x"BABBBBBB", x"C1C2C7CC", x"CECED0D3", x"D3D8DDDE", x"E0E5EAEB", x"EBEEEEEC", x"EBEBEAE8",
									 -- x"E7E6E6E6", x"E6E5E3E0", x"D9D5D1CE", x"CECFCFCF", x"D0CDCBCC", x"CFD1CFCD", x"D0D0D1D3", x"D6D9DADA",
									 -- x"DDDEE3EA", x"EEEFEEEF", x"EFEFEDEC", x"EBEBEBEC", x"EBEDEFEF", x"EDECECED", x"EBEDEEED", x"ECEAE7E4",
									 -- x"E1DFDCDA", x"D9D8D7D6", x"D7D6D4D4", x"D3D2D0CE", x"CFCCCBCD", x"CDCBCAC9", x"C3BFBCBA", x"BBBDBDBC",
									 -- x"BCBCBDBF", x"BEBCBCBE", x"BBBCB9B5", x"B4B6B7B5", x"B4B6B7B5", x"B3B2B1AF", x"B0B4B8B8", x"B5B2B1B0",
									 -- x"AEADABA9", x"A8A7A6A6", x"A3A4A4A2", x"A1A1A09E", x"9B9A9693", x"9597928A", x"8685827C", x"78777A7D",
									 -- x"89959696", x"9E9F9CA1", x"9B939090", x"8D8B8984", x"7F7C7B7E", x"858E9088", x"8678777E", x"7D7D7E7A",
									 -- x"75787770", x"69656464", x"65646361", x"5E61625D", x"5F5E5E5D", x"5D5C5C5C", x"5A5A5A5B", x"5C5D5B5A",
									 -- x"5F626164", x"5F585C5C", x"5A575657", x"56535354", x"57555354", x"54545658", x"57575859", x"5C5E5E5E",
									 -- x"5E636766", x"64656666", x"686A6B6C", x"6F75787A", x"81808183", x"82808287", x"858C8E8B", x"8B90928F",
									 -- x"8D898687", x"888B8F93", x"91939395", x"9B9C9B9D", x"A1A2A3A3", x"A4A5A7A8", x"A9ABABAB", x"ACAFB1B1",
									 -- x"B4B7BABB", x"BCBEC0C1", x"C3C7C9C8", x"C9CCCDCB", x"CECDCED1", x"D1CFCFD0", x"CDCECECC", x"CBCBCBCA",
									 -- x"C6C9C9C7", x"C7C8C8C6", x"CACACAC9", x"CACCCAC7", x"C7C4C2C1", x"BEB8B3B1", x"ADA7A19F", x"99908A88",
									 -- x"625E5C5D", x"5B595B5F", x"57565553", x"52504E4D", x"504C4C4B", x"48494A48", x"48464648", x"48484747",
									 -- x"44454747", x"46444444", x"47454445", x"45444548", x"46464646", x"4A4D4D4B", x"4E4C4A4A", x"4B4D4D4D",
									 -- x"4C4C4C4C", x"4F525454", x"52525455", x"53504F51", x"54535355", x"5758595B", x"5D626463", x"666B6B66",
									 -- x"6A6A6B6E", x"71747779", x"857F7C80", x"8384868A", x"8B8A8A8B", x"8F939597", x"95969799", x"99989695",
									 -- x"98959597", x"958F8E90", x"93959899", x"98989899", x"99969596", x"96959495", x"939B9E9F", x"A2A5A8AC",
									 -- x"ADACADB1", x"B5B9BFC5", x"C9C9CACC", x"CFD1D2D2", x"D3D5D6D9", x"DCDFDFDE", x"D9D5D2D1", x"CEC9C7C8",
									 -- x"C9C5C3C5", x"C4C1BCBA", x"B8BABAB7", x"B5B5B6B6", x"B7B4B1B1", x"B4B7B7B6", x"B6B6B6B6", x"B6B5B5B5",
									 -- x"B2B2B1B4", x"BABBB9BC", x"C0C2C5C9", x"CBCDD1D6", x"D6D7D8D9", x"DCDFE4E6", x"E6EAEDED", x"E9E6E6E6",
									 -- x"E8E6E4E3", x"E4E4E3E1", x"DBD6D2D1", x"D1D0D0D1", x"D3CFCBCA", x"CCCDCBC9", x"CACDCFCF", x"CFD3D6D7",
									 -- x"D8D9DCE3", x"EBF0EFED", x"EFEBE8E8", x"EAEDEEED", x"EEECECEE", x"EFEDECED", x"F1F0F0EF", x"EEECE9E7",
									 -- x"E6E2E0E0", x"DEDBDCE0", x"DBDAD8D5", x"D2D1D1D1", x"D2CCC8C7", x"C8C8C7C7", x"C1BDB9B8", x"BBBDBDBC",
									 -- x"BBBBBBBB", x"BABBBCBD", x"B5B7B6B3", x"B4B8B7B2", x"B3B3B1AE", x"ACADAFB1", x"AFB0B3B7", x"B6B1ADAB",
									 -- x"ABAAAAA9", x"A7A4A3A3", x"A3A3A2A0", x"9E9C9C9C", x"96939499", x"98908C8C", x"83857D7E", x"7A81828C",
									 -- x"91989D9D", x"9C9C9E9F", x"9C97908C", x"8D8E8A85", x"7A7E7F83", x"8D93918F", x"86837D79", x"797A7875",
									 -- x"74747370", x"6B676565", x"63646360", x"5E5E5D5B", x"5C5D5B59", x"585A5C5C", x"57585A5A", x"5A5B5C5E",
									 -- x"5B5B5B5A", x"5A5A5A5B", x"58515558", x"53535653", x"55545453", x"52535455", x"55585958", x"585A5D5E",
									 -- x"5E606263", x"63646667", x"68676B6C", x"6C707676", x"757C7C7D", x"817F808B", x"85878888", x"8B8C8A87",
									 -- x"8A888687", x"898B8B8A", x"8E8F8F92", x"9796979C", x"9F9F9FA2", x"A4A6A6A6", x"A9ABABA9", x"ABB1B3B0",
									 -- x"B2B5B9BC", x"BCBBBBBD", x"C1C3C5C5", x"C5C4C4C4", x"CDCBCCCF", x"CECBCACA", x"C9C8C7C7", x"C8C7C6C4",
									 -- x"C7C4C1C2", x"C4C6C4C3", x"CBC7C5C8", x"CBCBC9C8", x"C0BFBEBC", x"B8B3ADA9", x"A6A29D9A", x"958E8B8A",
									 -- x"5B5A5959", x"58565657", x"56545250", x"4F4E4D4D", x"4E4A4A4A", x"48484844", x"46464645", x"45454645",
									 -- x"46464645", x"42403E3D", x"43414041", x"41404244", x"44454545", x"47494947", x"4C4B4A49", x"49494949",
									 -- x"48494A4A", x"4A4C4E50", x"4F4F5152", x"504E4E50", x"54535354", x"55565759", x"5C5C5F62", x"63636567",
									 -- x"6768696C", x"6E727476", x"7E7B7C80", x"8383858A", x"8B8D8E8F", x"90929598", x"9797999B", x"9C9C9D9E",
									 -- x"9E9D9E9F", x"9B969699", x"96989B9D", x"9E9F9F9F", x"A19E9B9B", x"9B9B9C9E", x"989D9FA0", x"A5A9AAAE",
									 -- x"B7B5B5B7", x"B9BABEC2", x"C7C7C7C9", x"CBCDD0D1", x"D2D2D4D8", x"DBDDDEDE", x"DFDAD6D4", x"D2CDCAC9",
									 -- x"CAC6C5C6", x"C6C4C0BF", x"BDBEBCB9", x"B8B9B9B7", x"B8B8B9B9", x"BABABABA", x"B6B5B5B5", x"B6B5B3B2",
									 -- x"B3B3B2B4", x"B9B9B8BC", x"BCBEC3C8", x"CBCED2D7", x"D7D8D8D9", x"DADDDFE2", x"E5E8EBEC", x"EAE8E7E7",
									 -- x"E4E2E0DF", x"E0E0DFDE", x"DBD7D3D2", x"D1CFCDCD", x"D0CECCC9", x"C7C6C5C5", x"C7CBCCCB", x"CACDD0D2",
									 -- x"D5D6D9E0", x"E7ECEEED", x"EBE8E5E5", x"E7EAEDEE", x"EEECECEE", x"EFEEEEF0", x"F1F0F0F0", x"EFEDEAE8",
									 -- x"E9E5E4E5", x"E3E0E2E6", x"E3E0DCD9", x"D7D5D4D2", x"D2CDC9C9", x"CAC9C7C6", x"C2BEB9B8", x"B9BBBBBA",
									 -- x"BABABABA", x"B9B8B7B6", x"B5B3B2B3", x"B4B3B2B2", x"B5B2AFAD", x"ADAEAEAE", x"AFAFB2B5", x"B5B1AEAD",
									 -- x"A8A7A7A6", x"A5A3A1A0", x"9FA0A1A0", x"9D999796", x"94929294", x"938F8C8D", x"87877D7F", x"808A8D97",
									 -- x"949BA0A1", x"9F9D9A98", x"96938F8D", x"8D8C8882", x"7E7F7E81", x"8C929393", x"8A867F79", x"77777572",
									 -- x"7171706D", x"68646261", x"6564625D", x"5B5A5855", x"595A5855", x"54565858", x"59575553", x"5356595C",
									 -- x"5B5B5A59", x"58575757", x"57525557", x"52525452", x"55545352", x"51525556", x"53565857", x"575A5C5E",
									 -- x"5B5D5F61", x"63646667", x"6465696C", x"6B6E7272", x"74767579", x"82807B7E", x"84858586", x"8A8D8B88",
									 -- x"8C898685", x"86898C8D", x"898B8C91", x"9899999D", x"9D9D9EA1", x"A4A6A7A7", x"A8ABABAA", x"ADB3B4B1",
									 -- x"B2B4B7BA", x"B9B8B9BB", x"C0C0C0C2", x"C3C3C2C2", x"C8C6C5C6", x"C6C5C6C9", x"CCC7C1BE", x"BEC0C3C5",
									 -- x"C3C2C0C0", x"C1C2C3C3", x"C4C2C4C7", x"C8C6C3C2", x"BEBDBBB8", x"B4AEA9A5", x"A09C9895", x"928E8B8A",
									 -- x"58595856", x"56565655", x"54524F4D", x"4C4C4C4C", x"49464849", x"49494844", x"43454542", x"41434443",
									 -- x"45454443", x"4342403F", x"3E3D3C3D", x"3D3D3D3F", x"40414242", x"43444544", x"46474746", x"45444444",
									 -- x"45474848", x"4747494C", x"4D4C4D4E", x"4D4C4D50", x"53525153", x"54545658", x"5C595C62", x"625E6169",
									 -- x"68696A6C", x"6F727576", x"7A7B7F83", x"8584878C", x"8C8F9293", x"92929597", x"97999A9A", x"9B9EA2A4",
									 -- x"A2A3A5A5", x"A19C9DA1", x"9D9EA0A2", x"A4A5A4A4", x"A4A2A0A0", x"A1A0A1A2", x"9B9F9FA0", x"A6AAABAD",
									 -- x"B7B7B8BB", x"BCBEC0C3", x"C7C8C8C9", x"CACCD1D4", x"D1D0D3D7", x"D9D9DCDF", x"DFDAD6D6", x"D6D3CFCD",
									 -- x"CCC9C7C7", x"C8C7C6C5", x"C3C2BFBD", x"BDBEBCB9", x"B8BBBDBD", x"BBBABBBD", x"BABAB9BA", x"BAB9B6B4",
									 -- x"B5B6B4B5", x"B8B7B7BC", x"B6B9BFC6", x"CACDD1D4", x"D6D6D6D6", x"D6D7DADB", x"E2E5E8EA", x"EAE9E8E7",
									 -- x"E5E2E0DF", x"DFDEDEDC", x"DAD7D4D4", x"D3D0CDCD", x"CBCCCBC9", x"C5C3C5C7", x"C4C7C9C7", x"C5C7CACD",
									 -- x"D1D2D5DA", x"E0E4E7E7", x"E4E2DFDE", x"E0E4E9EC", x"EDEBEBEC", x"EDEEEFF1", x"F1F1F0F0", x"EFEEECEA",
									 -- x"ECE9E8E9", x"E8E7E8EC", x"EBE6E1DD", x"DBD9D6D3", x"D2CECACB", x"CCCAC7C6", x"C2BDB9B7", x"B8BABAB9",
									 -- x"B9B9B9B7", x"B6B3B1B0", x"B4B0AFB2", x"B2AFAFB2", x"B5B0ACAB", x"AEAFAEAC", x"B0B0B1B3", x"B2B0ADAD",
									 -- x"A8A8A7A6", x"A4A2A09E", x"9C9D9C9B", x"99969492", x"93939292", x"92919191", x"8F8D8587", x"8B94959A",
									 -- x"999DA1A1", x"9F9C9793", x"94939190", x"8F8C8680", x"7F818083", x"8C919090", x"85827C77", x"75757370",
									 -- x"71706F6C", x"68646260", x"61605D5A", x"5A5A5856", x"58595754", x"53545656", x"56565554", x"55555554",
									 -- x"58575655", x"54535352", x"53515354", x"504F5150", x"5252514F", x"4F515355", x"51545655", x"56595B5C",
									 -- x"5A5B5C5F", x"61626261", x"62626669", x"686A6F6F", x"6E74777A", x"7D7A797E", x"83828283", x"878A8986",
									 -- x"8787898A", x"8B8C8C8B", x"87898A8F", x"97999A9E", x"9C9C9EA1", x"A4A5A6A6", x"A7A9AAAA", x"ACB0B1AF",
									 -- x"B1B1B3B5", x"B4B4B5B8", x"BDBCBBBC", x"BFC0C0BF", x"C2C0BFBF", x"BFBFC0C2", x"C1C0BFBE", x"BFC1C2C2",
									 -- x"C1C0BFBE", x"BEBFC2C3", x"C2C3C4C4", x"C2BEBCBB", x"B9B8B5B2", x"AEA9A4A1", x"9C989493", x"918D8A88",
									 -- x"57585753", x"54575856", x"514F4D4B", x"4B4B4B4A", x"49474949", x"46464642", x"3F434340", x"3F424341",
									 -- x"43424142", x"44444443", x"3C3B3B3B", x"3C3B3C3C", x"3B3E3F3F", x"40424342", x"3F424444", x"41404042",
									 -- x"43444546", x"4646484B", x"4C4B4C4C", x"4C4B4C4F", x"51504F51", x"52535558", x"5A585A61", x"615D6067",
									 -- x"67686A6C", x"70737577", x"7B7C8085", x"8787898D", x"8E919495", x"94949495", x"999B9C9B", x"9C9FA4A6",
									 -- x"A5A6A8AA", x"A8A4A3A5", x"A5A4A3A4", x"A6A7A6A5", x"A4A3A4A6", x"A6A3A1A1", x"9FA3A2A2", x"A6AAABAD",
									 -- x"B3B6BABE", x"C0C2C4C5", x"C8CACACA", x"CACCD0D4", x"D1D0D2D6", x"D7D7DAE0", x"DFDCDBDA", x"DAD7D3D1",
									 -- x"CDCBC9C9", x"C9CAC9C9", x"C6C6C3C1", x"C0C0BFBD", x"BDBEBEBC", x"BABABCBF", x"BFC0C1C1", x"BFBDBBB9",
									 -- x"B7B9B7B6", x"B7B5B6BC", x"B7B9BEC5", x"C9CBCFD2", x"D5D5D4D3", x"D3D5D7D9", x"DEE0E3E6", x"E8E9E8E8",
									 -- x"E7E5E3E0", x"DFDEDDDD", x"DAD7D6D6", x"D6D4D2D1", x"CCCDCDCA", x"C7C5C6C8", x"C3C6C8C7", x"C4C5C8CC",
									 -- x"CDCFD3D6", x"D8DADCDD", x"DCDBD9D7", x"D7DCE2E6", x"ECEBEBEB", x"ECEDEEF0", x"F2F1F0EF", x"EFEFEEED",
									 -- x"EDEBEBEC", x"EBEAEBEE", x"EDE9E4DF", x"DCD9D5D3", x"D1CDCBCC", x"CDCBC9C7", x"C0BDB9B7", x"B8B9B9B9",
									 -- x"B9B8B5B3", x"B1B0AFAE", x"B1AEADAF", x"AFADAEB1", x"AFACA9AA", x"ADAFAEAC", x"B1B1B1B0", x"AFADABAB",
									 -- x"A8A8A7A5", x"A2A09D9B", x"9B999796", x"96969595", x"92949594", x"94949492", x"92949193", x"999B9797",
									 -- x"9C9D9E9E", x"9D9B9693", x"93949391", x"8F8C857F", x"7E828488", x"8F8E8886", x"7D7B7774", x"7474706C",
									 -- x"70706F6C", x"69666361", x"5E5C5A59", x"5A5A5958", x"57585855", x"54555555", x"53545555", x"54535251",
									 -- x"54545453", x"53525151", x"504F5050", x"4D4C4E4F", x"4E4E4E4D", x"4D4E5052", x"51535453", x"5457595A",
									 -- x"5A5A5A5C", x"5D5E5C5A", x"625F6164", x"63666D6F", x"6D727778", x"77777A80", x"807E7E80", x"83858481",
									 -- x"8083878B", x"8C8C8B8B", x"8A8B8A8B", x"9195999F", x"9D9EA0A1", x"A3A3A3A3", x"A6A8A8A7", x"A8ABABAA",
									 -- x"AEADAEAF", x"AFAFB1B4", x"B9B8B8B8", x"BABCBDBD", x"BDBDBDBE", x"BDBCBBBB", x"B9BBBEC0", x"C1C0BEBC",
									 -- x"BFBEBCBC", x"BDBFC1C2", x"C0BFBEBD", x"BBBAB9B9", x"B2B1AFAC", x"A9A6A2A0", x"9B989593", x"918C8783",
									 -- x"54565552", x"53555552", x"4F4E4C4B", x"4B4A4A49", x"4B494A48", x"423F403E", x"3D404140", x"4041413F",
									 -- x"41403E3F", x"40403F3D", x"3C3C3C3C", x"3C3C3C3B", x"3A3C3E3D", x"3E404141", x"3D404443", x"413F3F41",
									 -- x"42404144", x"46464749", x"4B4B4C4C", x"4B4A4C4E", x"504E4E50", x"51515356", x"5657595B", x"5E5F6060",
									 -- x"62646669", x"6D717375", x"7C7D7F83", x"8688898B", x"8F919395", x"97969594", x"9A9D9F9E", x"A0A3A6A7",
									 -- x"A9AAACAF", x"AFADAAA9", x"ACAAA7A7", x"A8A9A9A9", x"A8A7A7A9", x"A9A6A3A3", x"A2A8A8A6", x"A7A9AAAE",
									 -- x"B3B7BDC1", x"C4C5C5C5", x"C7C9CACA", x"C9CACCCF", x"D1D0D2D5", x"D6D6D9DE", x"E3E4E4E2", x"DED9D5D2",
									 -- x"CFCECCCA", x"CBCBCBCA", x"C6C8C7C4", x"C2C2C2C2", x"C3C2C1C0", x"BFBFC0C0", x"C0C3C5C5", x"C1BEBCBD",
									 -- x"B9BBBAB8", x"B7B5B5BB", x"BBBCBFC5", x"C9CBCED1", x"D5D5D3D2", x"D1D3D5D7", x"D9DBDEE1", x"E4E7E8E8",
									 -- x"E6E5E3E1", x"E0DFDEDE", x"DCD9D7D8", x"D8D7D6D6", x"D3D2D0CD", x"C9C7C5C5", x"C6C8CAC9", x"C6C4C7CA",
									 -- x"CBCED1D4", x"D4D4D5D5", x"D6D5D4D2", x"D1D5DBDF", x"E9EBECEC", x"ECEDEEEF", x"F2F0EEED", x"EEEFF0F0",
									 -- x"EEEDEDED", x"ECEBECED", x"ECE9E5E0", x"DAD6D4D3", x"D0CCCACC", x"CDCCCAC9", x"C1BEBAB9", x"B9B9B8B7",
									 -- x"B8B5B1AF", x"AEAEAEAF", x"AAABAAAA", x"AAABADAD", x"A9A9AAAB", x"ACADADAC", x"B1B1B0AE", x"ACABA9A8",
									 -- x"A5A6A5A1", x"9F9E9C99", x"9A989696", x"97979695", x"92969897", x"9695928F", x"94999B9B", x"A19F9B98",
									 -- x"9D9C9C9D", x"9D9A9592", x"90908F8D", x"8D8B8681", x"7E82868B", x"908C8380", x"7E7B7672", x"71726F6B",
									 -- x"6E6E6C6A", x"68656261", x"615E5B59", x"58565554", x"52545554", x"53535351", x"5353524F", x"4C4D5053",
									 -- x"53535353", x"52515050", x"4E4F4E4B", x"4B4B4C4F", x"4A4B4C4C", x"4C4D4D4E", x"50515251", x"52555656",
									 -- x"58575859", x"5B5C5B59", x"605C5F62", x"61646B6E", x"6E6D6E72", x"75787876", x"7B7B7C7F", x"8182807F",
									 -- x"81818182", x"84878B8E", x"898D8D8C", x"8F92969D", x"9E9FA1A2", x"A2A2A2A2", x"A5A6A5A4", x"A4A6A7A7",
									 -- x"AAA9A9AB", x"ABACAEB1", x"B4B5B5B5", x"B4B6B9BC", x"BABABBBB", x"BABAB9B7", x"BCBBBAB9", x"B8B7B7B7",
									 -- x"BCBAB7B8", x"BABDBDBD", x"B7B6B5B4", x"B6B7B7B6", x"ADACAAA8", x"A5A3A09E", x"99989592", x"8F8A837E",
									 -- x"53545555", x"5555514D", x"4F4E4C4B", x"4A4A4948", x"48464745", x"3F3E403F", x"3D3D3E40", x"40403E3D",
									 -- x"3D3D3C3C", x"3D3C3B3A", x"3C3D3D3C", x"3C3C3B39", x"3B3C3C3B", x"3C3E3E3E", x"3D404343", x"403E3E3F",
									 -- x"3F3D3D41", x"43434345", x"49494A4C", x"4B494A4C", x"4D4C4D4E", x"50505153", x"55585958", x"5B61615E",
									 -- x"60616468", x"6C707374", x"7E7E8084", x"878A8B8C", x"90919396", x"98999896", x"9A9D9F9F", x"A2A6A8A6",
									 -- x"ACACADB0", x"B2B2AFAC", x"B1AFADAC", x"ACADAEAF", x"AEABA9A9", x"A8A7A6A7", x"A4AAAAA7", x"A8A8A9AE",
									 -- x"AFB4BBBF", x"C3C6C7C6", x"C8C9CBCB", x"CBCBCCCD", x"D1D1D2D4", x"D6D8DBDD", x"E3E5E7E4", x"DFDBD8D6",
									 -- x"D2D2D0CF", x"CECFCECC", x"C8CACAC7", x"C5C5C6C6", x"C4C4C4C5", x"C6C5C3C1", x"C2C5C8C7", x"C4C0BFBF",
									 -- x"BCBDBBB9", x"B9B6B5BA", x"BABABDC2", x"C6C8CBCE", x"D1D1D0CE", x"CECED0D1", x"D4D6D9DC", x"DFE3E6E8",
									 -- x"E6E5E5E4", x"E3E2E2E1", x"DFDDDBDB", x"DBDAD9D9", x"D7D5D2CF", x"CECCCAC8", x"CDCDCDCC", x"C9C6C5C7",
									 -- x"CACDD0D2", x"D3D3D2D2", x"D3D2D1D0", x"CFD1D5D8", x"E3E7EBEC", x"EDEEEEEE", x"F0EEEDED", x"EEEFF0F1",
									 -- x"EEEFEFEF", x"EEEDEDED", x"EAE9E5DF", x"D9D5D3D3", x"CDCAC9CC", x"CECDCAC8", x"C2C0BDBA", x"B9B7B4B2",
									 -- x"B5B2AEAC", x"ABACADAC", x"A4A6A7A5", x"A5A7A8A8", x"A6A9ACAD", x"ADACABAC", x"AEAEAEAC", x"ABAAA8A7",
									 -- x"A2A4A3A0", x"9F9F9E9B", x"9A99989A", x"9B9A9592", x"97999C9D", x"9A969291", x"9BA0A29C", x"9F9C9A98",
									 -- x"9C9B9B9D", x"9D98918D", x"8D8C8A89", x"8B8B8884", x"81838487", x"8B878180", x"7E7A736F", x"70737473",
									 -- x"6E6D6B69", x"67646260", x"5E5C5957", x"55535253", x"50525352", x"51525250", x"5051514F", x"4D4C4E4F",
									 -- x"4F4F4F4F", x"4E4C4B4A", x"4E504B48", x"4A4B4A4D", x"484A4B4C", x"4C4B4B4B", x"4E4F4F4E", x"4F525352",
									 -- x"53545557", x"5A5C5C5D", x"5C5A5E63", x"6263676A", x"68696F73", x"72747572", x"77787B7F", x"81808081",
									 -- x"81818283", x"85888A8B", x"868C8E8E", x"91939599", x"9B9DA0A1", x"A2A2A2A2", x"A3A4A3A2", x"A2A3A5A7",
									 -- x"A7A6A6A8", x"A9A9ABAD", x"AEB0B2B1", x"AFB0B4B8", x"B5B6B5B4", x"B4B6B6B6", x"B8B8B7B6", x"B5B4B5B6",
									 -- x"B6B3B1B3", x"B6B8B7B5", x"B3B3B2B2", x"B2B2AFAB", x"AAA8A6A4", x"A19E9B99", x"9494938F", x"8A86807B",
									 -- x"55535355", x"56555251", x"4F4E4B49", x"49484848", x"46434344", x"42434441", x"403C3B3E", x"403D3B3B",
									 -- x"393A3B3C", x"3B3B3B3B", x"3A3C3D3B", x"3A3A3936", x"3A3A3938", x"393C3D3B", x"3B3D3F40", x"3E3C3C3D",
									 -- x"3E3C3D40", x"403D3E41", x"4344474A", x"49474748", x"4848494D", x"4E4F5052", x"55585856", x"585E615F",
									 -- x"6163666A", x"6E717475", x"7B7E8285", x"888B8E90", x"91939598", x"9A9B9C9C", x"9B9E9FA0", x"A4A9A9A6",
									 -- x"ACADAEAF", x"B1B2B1B0", x"B4B3B3B2", x"B1B1B2B3", x"B1AEABAA", x"A9A9A9AB", x"A7ACACAA", x"ACACACAF",
									 -- x"ADB2B8BC", x"C1C7CACA", x"CBCCCDCE", x"CECFCFCF", x"D2D5D6D6", x"D9DFE1DF", x"E2E4E4E1", x"DEDEDCDA",
									 -- x"D5D6D6D4", x"D3D4D2CF", x"CCCDCCC9", x"C8C9C9C9", x"C5C5C6C8", x"C9C9C7C5", x"C6C7C8C8", x"C7C5C2C0",
									 -- x"BEBFBCBB", x"BBB7B5B9", x"B9B9BCC1", x"C5C6C7C9", x"CACBCCCD", x"CCCCCCCC", x"CFD2D5D8", x"DBDEE4E7",
									 -- x"E8E9E9E8", x"E7E5E5E4", x"E3E1E0E1", x"E1DFDDDD", x"DAD9D7D6", x"D5D4D2D1", x"D3D2D1D1", x"CECAC7C7",
									 -- x"CBCCCED0", x"D1D1D1D0", x"CFCFCFCE", x"CECFD1D2", x"D8DFE6EA", x"ECEEEEEC", x"ECECECED", x"EFEFEFEF",
									 -- x"EDEEEFEF", x"EEEDEDED", x"EAE7E2DD", x"D8D4D1D0", x"CAC9C9CD", x"CFCDC8C6", x"C2C0BEBB", x"B8B5B1AF",
									 -- x"B0AEACAB", x"ABAAA8A6", x"A3A2A3A5", x"A4A2A2A5", x"A4A8ACAF", x"AFAEACAC", x"ACADADAB", x"A9A9A6A3",
									 -- x"A2A4A3A0", x"9FA1A19E", x"9B9A999B", x"9C9B9590", x"99999C9E", x"9C979698", x"9FA1A096", x"9A979896",
									 -- x"99989899", x"97928C89", x"8A888685", x"888B8883", x"83828080", x"83807C7D", x"79756F6C", x"6E737575",
									 -- x"6E6C6966", x"64615F5D", x"5A585756", x"54515356", x"52535350", x"50515151", x"4D4D4E4F", x"504E4B48",
									 -- x"4A4A4A4A", x"49484746", x"4B4E4844", x"49494546", x"46474849", x"48484848", x"4A4B4B4B", x"4C4F504F",
									 -- x"50515354", x"5557595B", x"5C595D62", x"61606466", x"62667173", x"6D707675", x"75777B7E", x"7E7D7F82",
									 -- x"7E808286", x"898A8987", x"878C8D8D", x"93959495", x"999B9EA0", x"A1A1A1A2", x"A2A2A2A2", x"A1A1A3A4",
									 -- x"A5A4A4A7", x"A8A7A7A9", x"AAABACAB", x"AAABAEB1", x"B0B1B1B0", x"B0B2B2B0", x"AFB1B4B6", x"B5B5B4B4",
									 -- x"AFAEAEB0", x"B2B2B1AF", x"B1B2B1AE", x"ACAAA8A4", x"A6A5A2A0", x"9D9A9694", x"9192908A", x"85817E7B",
									 -- x"57514F51", x"53535457", x"504E4A48", x"47474848", x"4B464445", x"4545443E", x"423B383D", x"3F3B3839",
									 -- x"393A3C3B", x"39373737", x"393B3B39", x"38383633", x"38373535", x"383C3D3B", x"36383B3C", x"3B3B3B3B",
									 -- x"3E3D3E40", x"3E3A3A3F", x"3F404447", x"47454546", x"4343464B", x"4E4F5153", x"53555553", x"53585D60",
									 -- x"6263666A", x"6E717375", x"757B8285", x"87898D90", x"9194989A", x"9B9C9FA1", x"A0A2A2A2", x"A7ACACA7",
									 -- x"ADAFAFAF", x"B0B1B4B5", x"B5B6B7B6", x"B4B3B3B4", x"B2B0AEAE", x"AEADACAD", x"ADB1B0AF", x"B2B4B2B3",
									 -- x"B1B6B9BC", x"C1C7CCCD", x"CDCDCDCE", x"CFD1D1D0", x"D4D8D9D8", x"DDE5E7E3", x"E8E8E5E0", x"DFDFDDDA",
									 -- x"D8DADAD9", x"D8D8D5D2", x"D0CFCDCB", x"CBCDCCC9", x"C8C8C9C9", x"CACBCCCD", x"C8C6C5C6", x"C8C7C3BF",
									 -- x"BFBFBDBC", x"BCB8B6B9", x"BCBCBFC4", x"C7C7C7C7", x"C7C9CDCF", x"CFCFCECD", x"CCCFD3D5", x"D7DCE2E7",
									 -- x"EBEBEBEA", x"E8E5E4E3", x"E5E4E4E6", x"E7E5E2E1", x"E1E1DFDD", x"DBD9D7D7", x"D6D4D4D5", x"D3CECAC9",
									 -- x"CBCBCCCD", x"CECFCECE", x"CBCCCCCD", x"CECECECE", x"CFD8E2E7", x"EAEDECEA", x"EAEAECEE", x"F0F0EFED",
									 -- x"ECEDEEEE", x"EDEDEDEC", x"EAE6DFDB", x"D7D4D0CD", x"C9C8CACE", x"D0CDC7C3", x"C0BFBDBB", x"B8B5B1AE",
									 -- x"ACABABAB", x"ABA8A4A0", x"A5A0A1A7", x"A59E9FA5", x"A3A7ACB0", x"B1B1AFAD", x"ACAEAEAB", x"A9A7A4A0",
									 -- x"A2A4A29E", x"9DA0A09D", x"9D9A9899", x"9B9A9692", x"9795989C", x"9B97999E", x"9A9B9A90", x"97959896",
									 -- x"98959392", x"908C8888", x"88858181", x"8587847E", x"82817C7C", x"7D797577", x"74726E6C", x"6D706F6C",
									 -- x"6C696561", x"5F5D5A58", x"5A595857", x"53505257", x"5353514E", x"4C4E5051", x"504C4747", x"4A4B4946",
									 -- x"4848494A", x"49494847", x"484C4541", x"47464040", x"45454545", x"45444546", x"47484948", x"4A4D4F4E",
									 -- x"50515251", x"51515355", x"5E5A5C60", x"5E5E6366", x"6462676B", x"6C747A75", x"75777A7C", x"7B797C81",
									 -- x"7E7D7D7F", x"84888989", x"8B8D8A8B", x"92969594", x"989A9D9F", x"9F9FA0A0", x"A2A2A2A2", x"A09F9FA0",
									 -- x"A4A3A4A7", x"A7A6A6A6", x"A8A7A7A7", x"A7A9ABAC", x"ACAFB1B0", x"B0B0ADA9", x"AEAFB0B0", x"AFAFB0B1",
									 -- x"AAACAEAF", x"B0AFADAC", x"AAADACA7", x"A4A4A5A5", x"A2A19F9E", x"9B979491", x"90918F87", x"817E7C7B",
									 -- x"55555756", x"51505251", x"4D4C4B4B", x"4C4C4A48", x"4D4D4D4B", x"4A494440", x"3F3E3D3C", x"3B3A3A39",
									 -- x"393B3D3D", x"3A373534", x"36373839", x"38363432", x"36373534", x"383D3C37", x"37383838", x"393A3734",
									 -- x"3B3A3A3B", x"3B3B3A39", x"3D414442", x"41434545", x"4646474A", x"4A494C4F", x"52515154", x"55575B60",
									 -- x"6263666C", x"72757574", x"7A7D8287", x"87878C93", x"9496999B", x"9C9EA1A4", x"A4A5A6A8", x"AAABACAC",
									 -- x"ACB1B0AE", x"B1B3B4B6", x"B5B3B1B1", x"B2B6B8BA", x"B4AFAEB2", x"B4B2AFB0", x"AFB4B8B9", x"B9BAB9B7",
									 -- x"B8B8BABE", x"C1C5CBD2", x"D0D1D2D2", x"D0D0D0D1", x"D4D7DADC", x"E1E6E8E7", x"E6E5E2DE", x"DDDEDEDC",
									 -- x"DADCE0E0", x"DEDCDADA", x"D8D5D3D2", x"D0CECDCF", x"CCCACBCD", x"CFCFCFD0", x"C7CCCBC8", x"C8C7C7C9",
									 -- x"C3C1BEBC", x"BCBCBBBB", x"BBC0C5C7", x"C7C7CBCE", x"CBCECFCE", x"CDCECECC", x"CBCCCDD1", x"D6DADDDE",
									 -- x"E7E7E8E9", x"E9EAEAEA", x"E5E6ECEF", x"ECEBEAE7", x"E6E6E6E4", x"E0DDDDDD", x"D7D7DBDC", x"D4CFCFCE",
									 -- x"CECDCCCC", x"CBCBCDD0", x"D1D0CFCE", x"CECFD0D1", x"D1D3D8E1", x"E7E8E8E9", x"E9ECEEEC", x"EDF0EFEB",
									 -- x"ECEEEFEE", x"ECEAE9E9", x"E8E3DFDD", x"D9D2CCC9", x"C2C6CCD0", x"D0CDC8C6", x"C6C0BBBA", x"B7B0ADAD",
									 -- x"AAABAAA8", x"A6A7A7A5", x"A3A3A29E", x"9C9D9E9D", x"9EA1A5A8", x"A9A9A9A9", x"AEB0AEA9", x"A7A7A4A0",
									 -- x"9F9F9F9B", x"9A9F9F97", x"97989998", x"96949292", x"91979B9A", x"9A9D9E9C", x"9D989693", x"8D8D9191",
									 -- x"92908D8C", x"8B8A8684", x"7B7D8080", x"7E818079", x"7E7D7A78", x"78757377", x"726E6B6B", x"6C6B6A6A",
									 -- x"6768645F", x"5F605D58", x"55555656", x"5654514F", x"524E4C4D", x"4E4D4C4B", x"4E4A4944", x"46464249",
									 -- x"45464848", x"45434549", x"45474846", x"43414243", x"41404749", x"41414644", x"45464848", x"4A4C4D4D",
									 -- x"4F4E4F51", x"52525251", x"56585A5D", x"5E5F5E5D", x"6563666D", x"71707173", x"78757579", x"7D7E7D7C",
									 -- x"7C7F8284", x"84858789", x"8F89888F", x"96969492", x"97999C9D", x"9B989A9F", x"9B9F9F9D", x"9B9D9FA0",
									 -- x"A49FA0A3", x"A4A6A6A1", x"9FA2A4A4", x"A3A2A3A5", x"A6A7A8A9", x"AAAAAAAA", x"ACABABAD", x"AEADAAA8",
									 -- x"AAABACAB", x"AAA9A9AA", x"A9A7A4A3", x"A5A6A29C", x"9C9B9C9C", x"9A969291", x"948D8887", x"85807C7B",
									 -- x"52505355", x"53545553", x"50515150", x"4D4C4C4D", x"4C4D4E4D", x"4D4A4540", x"41403E3C", x"3A3A3A3A",
									 -- x"38393A3A", x"39373636", x"33343536", x"36363434", x"34353331", x"34383834", x"35373838", x"38393735",
									 -- x"3B3B3A3A", x"3A3A3A3A", x"3A3D3F3F", x"4042413F", x"42424447", x"4848494C", x"4D4D5054", x"56585C60",
									 -- x"6465676C", x"70747778", x"7D7F8386", x"888A8F96", x"95989C9F", x"9FA0A1A3", x"A4A6A9AC", x"AEAEAEAE",
									 -- x"AEB2B0AE", x"B0B2B2B4", x"B6B6B6B7", x"B8B8B8B7", x"B5B1B0B4", x"B7B5B4B5", x"B3B7BBBC", x"BCBEBEBC",
									 -- x"BDBDBFC2", x"C3C6CCD3", x"D3D3D2CF", x"CDCDCECF", x"D3D7DBDC", x"DEE3E7E9", x"E5E4E2DF", x"DFE0DFDD",
									 -- x"DBDCDDE0", x"E2E2E1E0", x"DDDAD7D6", x"D5D2D2D3", x"D2D1D0D2", x"D3D2D1D1", x"CDD1CFCB", x"CBCBC9CB",
									 -- x"C8C6C3C2", x"C2C2C1C0", x"BEC1C4C7", x"C9CBCDCE", x"CACDCECE", x"CED0D0CF", x"CECFD1D3", x"D5D7DADC",
									 -- x"E0E1E4E7", x"E9EAEAEA", x"E8E9EFF2", x"F0EFF0ED", x"EEEDEBE8", x"E6E2DFDE", x"DBDADFE2", x"DCD6D3CF",
									 -- x"D1CFCDCC", x"CCCCCED0", x"CECECFD0", x"D1D1D1D1", x"D2D2D5DC", x"E0E1E2E3", x"E6EAECEB", x"ECEEEDE9",
									 -- x"EDEEEFEE", x"ECEAEAEA", x"E7E2DDDB", x"D9D3CDCA", x"C5C9CED1", x"D1CDC9C6", x"C0BEB9B5", x"B3B2B0AE",
									 -- x"A9AAA8A5", x"A3A3A2A0", x"A19F9D9B", x"99999A9B", x"9E9F9FA0", x"A2A5A8AB", x"ACAFAEA9", x"A5A5A29F",
									 -- x"A09FA09E", x"9C9E9D95", x"98979594", x"92908E8C", x"8E949797", x"989B9C9A", x"9B979592", x"8C8C8E8D",
									 -- x"8E8C8A88", x"87858280", x"7B7C7E7D", x"7B7D7E78", x"79797776", x"77737073", x"6F6C6969", x"6A686767",
									 -- x"6663605E", x"5D5B5958", x"52525354", x"5453504F", x"4D4D4B49", x"4A4C4A46", x"47444442", x"46463F44",
									 -- x"45444445", x"44434445", x"42444443", x"41404143", x"42404345", x"40424744", x"47484949", x"494C4C4B",
									 -- x"4B4D4F51", x"5251504F", x"54585B5A", x"5A5B5C5C", x"6362656A", x"6C6B6E73", x"7475787A", x"7A787A7D",
									 -- x"7B7D8081", x"81838588", x"8B88878A", x"8F929496", x"9696989A", x"99969597", x"9C9C9C9C", x"98959598",
									 -- x"A09C9EA0", x"A1A3A39F", x"9E9E9D9D", x"9D9FA1A3", x"A2A3A5A6", x"A6A6A5A5", x"A5A4A4A5", x"A7A8A7A6",
									 -- x"A4A6A8A8", x"A7A5A5A5", x"A6A5A3A1", x"A1A19D97", x"9A989695", x"93908F8F", x"8B878484", x"827D7A7B",
									 -- x"53505254", x"53535350", x"54535150", x"4F4E4D4D", x"4B4D4F4E", x"4E4B4540", x"413F3E3D", x"3C3C3C3C",
									 -- x"3A393938", x"38373635", x"35353534", x"33323131", x"30323231", x"33363532", x"32343636", x"37383837",
									 -- x"3A3A3939", x"3838393A", x"393B3C3E", x"41423F3C", x"3E3E4043", x"4545474A", x"494C5055", x"58595B5E",
									 -- x"6365676A", x"6D71767A", x"7E808388", x"8B8E9296", x"969A9FA2", x"A3A2A3A3", x"A7A9ADB0", x"B2B2B1B0",
									 -- x"B1B4B3B0", x"B2B3B3B6", x"B6B7B7B8", x"B9B8B7B6", x"B9B5B4B7", x"BABAB9BB", x"B9BCBEBF", x"C0C2C3C2",
									 -- x"C4C5C7C8", x"C8C9CED3", x"D5D3D1CE", x"CBCCCED1", x"D0D5D8D8", x"D9DEE4E8", x"E6E6E4E2", x"E1E1DFDD",
									 -- x"DCDADADD", x"E3E7E7E6", x"E3E0DEDD", x"DBD9D9DA", x"D9D7D5D6", x"D5D3D1D0", x"D0D3D0CD", x"D0D0CDCE",
									 -- x"CBCAC8C7", x"C7C6C5C4", x"C4C4C6C9", x"CDD0D0CF", x"CDCFD0D0", x"D1D2D2D1", x"CCCED0D1", x"D2D4D7DA",
									 -- x"D8DBE0E4", x"E8E9E9E9", x"E8E9EEF3", x"F2F4F6F4", x"F4F2EFED", x"EBE8E4E0", x"E1DEE2E5", x"E2DDD9D4",
									 -- x"D4D1CECE", x"CECFD0D3", x"CFD0D1D3", x"D4D5D5D4", x"D5D4D4D7", x"D8D9D9DA", x"E3E8EBEB", x"EDEFEDEA",
									 -- x"EBEBEBEB", x"E9E8E8E8", x"E5E1DCDB", x"D9D6D1CE", x"CBCED1D3", x"D2CDC9C6", x"BDBDB9B2", x"B1B3B2AE",
									 -- x"AAAAA9A5", x"A3A2A19F", x"9F9B9998", x"9694969A", x"9D9C9C9C", x"9EA3A8AC", x"A9ACACA7", x"A3A2A19F",
									 -- x"A09D9D9E", x"9B9B9B97", x"97959291", x"9191908E", x"8E929698", x"9A9D9C99", x"96939290", x"8A898A88",
									 -- x"89888785", x"82807E7D", x"78787977", x"74777873", x"73747271", x"726D6A6C", x"6B696768", x"68666667",
									 -- x"635E5B5C", x"5A555458", x"51515151", x"514F4D4C", x"494B4945", x"464A4842", x"423F403F", x"43443D41",
									 -- x"44403E40", x"42424140", x"4141413F", x"3D3D3E40", x"423F3F40", x"3F424644", x"45464646", x"46484948",
									 -- x"4A4C4E4F", x"4F4F4F50", x"51575A56", x"55585B5B", x"60616467", x"66666B72", x"71737678", x"7776787B",
									 -- x"7C7D7E7F", x"80818486", x"8A8B8A88", x"898C9092", x"93929395", x"95929090", x"97949599", x"98939399",
									 -- x"99979A9C", x"9B9D9E9B", x"9C9A9897", x"999B9D9D", x"9C9D9FA1", x"A1A19F9E", x"A09F9E9E", x"A0A3A3A2",
									 -- x"9FA1A2A2", x"A1A0A0A0", x"A0A09F9D", x"9C9B9894", x"98969392", x"908D8C8D", x"8A878584", x"7F787678",
									 -- x"53505152", x"5050514E", x"55504C4B", x"4E4E4B48", x"4B4D4E4D", x"4D4A4540", x"3D3D3E3F", x"40403F3E",
									 -- x"3C3A3939", x"3A3A3837", x"35353534", x"3331302F", x"292D2F30", x"30323230", x"2E313435", x"36383A3A",
									 -- x"39383737", x"38393838", x"3A3A3C3E", x"40403D3B", x"3C3C3D3F", x"41444749", x"4A4D5256", x"58595A5C",
									 -- x"61646769", x"6A6F757B", x"7D80868C", x"91939495", x"999CA1A4", x"A4A4A5A6", x"AAACAFB2", x"B4B5B5B4",
									 -- x"B5B8B6B5", x"B8B8B8BB", x"BAB9B7B7", x"B8B9BBBB", x"BDBAB8BA", x"BCBCBDBE", x"BEBFC1C2", x"C4C5C5C5",
									 -- x"C7CACDCE", x"CDCDCFD2", x"D3D2D0CE", x"CCCED1D4", x"CFD2D4D5", x"D7DCE3E8", x"E9EAE9E6", x"E4E2E0DD",
									 -- x"DCDAD8DA", x"DFE4E7E7", x"E8E6E4E3", x"E2E1E1E2", x"E0DCD9D8", x"D7D4D2D1", x"D0D2D0CE", x"D3D4D2D2",
									 -- x"CECECDCC", x"CAC9C7C6", x"CAC9CACD", x"D1D3D3D1", x"D2D3D5D6", x"D6D6D3D1", x"CECFCFD0", x"D2D4D6D8",
									 -- x"D6D8DCE0", x"E3E4E4E4", x"E3E3E9EE", x"EFF3F6F5", x"F2F2F2F0", x"EFEDE9E5", x"E6E1E2E4", x"E1DFDFDC",
									 -- x"D8D5D2D3", x"D3D3D4D5", x"D5D5D5D6", x"D7D8DADB", x"D9D8D7D6", x"D5D5D4D5", x"DFE4E8EA", x"ECEEEEEC",
									 -- x"EAEAE9E9", x"E8E7E7E7", x"E1DFDDDA", x"D8D6D4D3", x"CFD1D4D4", x"D2CDC8C6", x"C0BEBAB4", x"B2B2B0AC",
									 -- x"ABAAA8A6", x"A3A2A1A0", x"9E999798", x"96929399", x"97999B9D", x"A0A3A7A9", x"A5A8A9A5", x"A1A0A09F",
									 -- x"9F999899", x"97979A99", x"96949291", x"90919192", x"8F929598", x"9C9D9A95", x"92908F8C", x"87878885",
									 -- x"86868583", x"7F7D7B7B", x"74747573", x"6F70716D", x"6E6E6C6B", x"6B676365", x"66646364", x"65646465",
									 -- x"5F5C5958", x"55515254", x"5150504F", x"4E4C4948", x"47484744", x"45474541", x"413F3F3C", x"3F403C42",
									 -- x"403D3B3D", x"40403E3E", x"41403F3D", x"3B3A3B3B", x"3F3D3D3D", x"3D3F4142", x"41424342", x"43464746",
									 -- x"4A4C4C4A", x"494B4F52", x"4F555753", x"52585C5C", x"5E606365", x"65656A70", x"72727276", x"7A7C7B7A",
									 -- x"7E7E7E7F", x"7F818486", x"898D8E8A", x"888B8C8C", x"8E8E8E8F", x"8F8E8D8D", x"8E8C8E93", x"95939599",
									 -- x"92929598", x"96979997", x"99989797", x"97979797", x"97989B9D", x"9D9D9C9B", x"9E9D9C9C", x"9D9FA09F",
									 -- x"9C9D9D9D", x"9C9C9EA0", x"98999A9A", x"99979593", x"95939291", x"8F8B8989", x"8B878482", x"7D777576",
									 -- x"4C4B4E4F", x"4C4E5252", x"504E4B4A", x"4B4B4A48", x"4B4C4C4C", x"4C4B4844", x"3F3E3D3E", x"40424241",
									 -- x"3B3A3A3C", x"3D3E3D3C", x"34353535", x"34333130", x"292A2B2A", x"2A2B2D2E", x"2D303333", x"34363939",
									 -- x"3A383638", x"3B3B3936", x"39393A3B", x"3B3B3A3A", x"3C3C3B3C", x"3F444749", x"4C4F5356", x"585A5C5D",
									 -- x"61656A6C", x"6D70777C", x"7F83898F", x"94989998", x"A0A3A5A6", x"A6A6A8AA", x"ABACAFB2", x"B5B7B9BA",
									 -- x"B9BCBBBA", x"BDBCBBBF", x"BFBDBBBA", x"BBBCBEC0", x"BEBCBBBC", x"BEBFC0C1", x"C1C1C3C5", x"C6C6C6C6",
									 -- x"C9CDD1D3", x"D3D3D2D2", x"D3D2D1CF", x"CECED0D2", x"D0D0D0D3", x"D8DDE3E7", x"EAECEBE8", x"E6E5E3E1",
									 -- x"DFDDDBDA", x"DCE0E4E7", x"EBEBEAE9", x"E9E9EAEA", x"E7E2DCDA", x"D9D7D6D6", x"D2D4D2D1", x"D7D9D6D5",
									 -- x"D3D3D2D0", x"CECCCACA", x"CBCCCFD1", x"D3D5D6D7", x"D9D9DBDD", x"DDDAD6D3", x"D5D3D1D2", x"D5D8D8D8",
									 -- x"D9DADBDC", x"DDDEDEDE", x"DFDEE3E7", x"E9EDF1F0", x"EEF1F4F2", x"F1EFEDEA", x"E7E3E3E4", x"E1E0E2E1",
									 -- x"DDDBDADA", x"D9D7D7D7", x"DADADADB", x"DBDCDDDD", x"DDDDDBD8", x"D6D4D3D3", x"DCE0E5E8", x"E9EAEAE9",
									 -- x"EAEAE9E9", x"E8E7E7E6", x"DFE0DEDA", x"D6D3D3D4", x"D1D3D5D5", x"D2CDC8C5", x"C4BFBBBA", x"B6B1ADAC",
									 -- x"A9A8A6A3", x"A19E9D9D", x"9B979698", x"96919196", x"93959A9D", x"A0A2A3A4", x"A5A8A9A6", x"A19F9F9F",
									 -- x"9E989797", x"95959898", x"94949391", x"8E8E9092", x"90909192", x"95969491", x"908E8D89", x"85878885",
									 -- x"83838280", x"7D7A7878", x"71717271", x"6C6C6C69", x"696A6766", x"66636063", x"62605F60", x"605F5F5F",
									 -- x"5B5C5954", x"5051514F", x"504F4D4C", x"4B494745", x"48444446", x"46434142", x"3F3F403C", x"3C3B383F",
									 -- x"3B3A3A3B", x"3C3C3C3E", x"403F3C3A", x"39393939", x"3A3C3C3B", x"3B3B3C3F", x"40414141", x"42454646",
									 -- x"484A4A47", x"474A4E50", x"4F535451", x"53595C5A", x"5C5D5F62", x"6466686B", x"6F6F7175", x"797D7D7D",
									 -- x"7D7E7E7E", x"7F818384", x"86898A88", x"888B8C8A", x"8A8B8B8A", x"88888A8B", x"8B8B8B8B", x"8D8F9090",
									 -- x"8F8F9394", x"92939594", x"95969695", x"93939495", x"94959799", x"9A9B9A99", x"9A9C9C9B", x"9C9E9D9B",
									 -- x"999A9B9C", x"9B9B9D9E", x"95969798", x"98959493", x"92908E8E", x"8B888686", x"85807D7D", x"7B787778",
									 -- x"49494C4C", x"494A4F50", x"4A4C4E4C", x"49484A4E", x"4A4B4B4A", x"4B4D4B48", x"44403C3B", x"3D404142",
									 -- x"3F3F3E3E", x"3D3D3B3A", x"38383837", x"3533302E", x"302F2B28", x"27292C2E", x"2D303130", x"31343536",
									 -- x"39383739", x"3C3C3936", x"3938393A", x"3938393A", x"3B3B3B3B", x"3E444748", x"4B4F5355", x"575B5E60",
									 -- x"62676D70", x"71747A7F", x"85888B8F", x"949A9E9F", x"A8A9AAA9", x"A8A8AAAC", x"AAABADB1", x"B4B8BCBE",
									 -- x"BCBFBEBE", x"C0BEBCC0", x"C0BFBEBE", x"BEBEBEBE", x"BEBDBDBE", x"C0C2C3C4", x"C3C3C4C7", x"C9C9C8C8",
									 -- x"CCD0D3D6", x"D8D9D7D5", x"D6D6D5D2", x"CFCDCDCD", x"CECDCED2", x"D7DCE1E5", x"E9EAEBE9", x"E8E8E8E8",
									 -- x"E5E5E2E0", x"DFE1E6EB", x"F0F1F1F1", x"F1F2F2F1", x"EBE4DEDC", x"DBDAD8D8", x"D7DAD8D7", x"DCDCD9D8",
									 -- x"D7D7D5D2", x"D0CECECE", x"CCCFD3D5", x"D7D9DCDF", x"E0DFE1E3", x"E3DFD9D6", x"D3D0CFD1", x"D6DBDCDB",
									 -- x"DCDCDAD9", x"D9D9DADA", x"DEDDDFE2", x"E3E6E9E7", x"EBF1F5F4", x"F3F3F2EF", x"E7E5E7E9", x"E6E4E3E1",
									 -- x"E2E1E1E1", x"DFDCDADB", x"DCDEE0E2", x"E2E1DEDD", x"DFE0DEDA", x"D7D6D5D4", x"DFE2E6E7", x"E7E6E5E5",
									 -- x"E8E7E6E6", x"E5E4E3E2", x"E2E3E2DC", x"D7D4D4D4", x"D1D3D5D5", x"D2CDC8C5", x"C5BFBCBC", x"B9B1ADAD",
									 -- x"AAA7A5A3", x"A09C9A9A", x"97949495", x"938F8F91", x"9496999C", x"9EA0A2A3", x"A7A8A8A5", x"A19E9D9D",
									 -- x"9C9A9A99", x"95959593", x"8F919291", x"8E8F9296", x"92908D8C", x"8D8F8F8E", x"8E8C8B88", x"84878883",
									 -- x"807F7E7B", x"79767473", x"706F706F", x"6A686967", x"65666363", x"64615F62", x"625F5D5E", x"5E5D5B5A",
									 -- x"58595750", x"4E504F4C", x"4B4A4948", x"47464544", x"46414145", x"45403E41", x"3B3B3F3C", x"3C393338",
									 -- x"3838383A", x"39383A3C", x"3C3A3838", x"39393938", x"363B3B3A", x"3B39383C", x"3E3F3F3E", x"3E414242",
									 -- x"43474847", x"474A4C4B", x"4F515252", x"54575856", x"59595B5E", x"62646464", x"63696F70", x"7073777B",
									 -- x"7A7A7B7C", x"7D7E7E7F", x"84858483", x"83868787", x"88898885", x"83838587", x"8A8A8886", x"888C8C8A",
									 -- x"8E8D9091", x"8F909291", x"91929190", x"8E8E9296", x"93939496", x"97979898", x"94979898", x"999B9B99",
									 -- x"94979A9C", x"9B9A9999", x"95959597", x"96939191", x"928F8B89", x"87848485", x"827D7B7C", x"7B777576",
									 -- x"4A494B4B", x"48484948", x"47494B4B", x"49494B4D", x"4A4A4A49", x"4A4B4946", x"44403C3A", x"3C3D3E3D",
									 -- x"42413F3D", x"3A383838", x"3A393837", x"35333130", x"3533302D", x"2C2C2D2E", x"2C2D2D2D", x"2F323333",
									 -- x"36363738", x"39383736", x"38363538", x"39393839", x"393A3A3B", x"3E444646", x"4B4F5355", x"575C6061",
									 -- x"62676D70", x"72757A7E", x"878A8D8F", x"939A9FA1", x"A8AAACAC", x"ABAAAAAB", x"ACADAEB1", x"B4B8BBBD",
									 -- x"BDC0C0C1", x"C3C0BEC2", x"C0BFBFBF", x"BFBFBFBE", x"C0C0C0C1", x"C2C4C5C6", x"C6C5C5C9", x"CBCCCCCE",
									 -- x"D1D3D5D8", x"DBDEDDD9", x"D8D9D8D5", x"D1CFCECE", x"CECDD0D4", x"D7DADFE4", x"E6E8E9E8", x"E8EBEDED",
									 -- x"ECEBE9E7", x"E6E8EEF2", x"F6F8F9F9", x"F9FBFAF8", x"ECE6E0DF", x"DEDCDAD9", x"DBDFDEDD", x"E0E0DBDA",
									 -- x"DCDBD8D5", x"D3D2D3D5", x"D3D5D9DB", x"DDE0E3E6", x"E8E6E6E7", x"E6E0DAD7", x"CFCECDD0", x"D5D9DCDD",
									 -- x"DDDBD9D7", x"D7D7D9DA", x"DDDBDDDF", x"DFE2E4E2", x"E8EEF3F4", x"F6F8F6F2", x"EBE7E9ED", x"EBE8E4DF",
									 -- x"E4E5E6E6", x"E3E0E1E4", x"E2E3E6E7", x"E7E5E3E1", x"E2E2E1DC", x"D9DADAD9", x"E1E4E6E7", x"E6E4E3E3",
									 -- x"E3E2E2E1", x"E1E0DDDB", x"E2E2E0DB", x"D8D7D5D3", x"D1D3D6D6", x"D3CEC9C6", x"C4C1BDBA", x"B7B2AEAC",
									 -- x"ABA8A5A4", x"A09C9A9B", x"94939391", x"8F8E8E8E", x"9697999B", x"9C9E9FA1", x"A4A4A3A2", x"9F9C9B9A",
									 -- x"9A9A9B97", x"9394948F", x"8D8F908F", x"8E8F9194", x"908E8D8C", x"8C8B8A89", x"8A898985", x"8284847E",
									 -- x"7E7C7A78", x"7674716F", x"6E6C6D6B", x"65646665", x"61626160", x"625E5B5E", x"5F5A5859", x"5C5B5755",
									 -- x"5554514E", x"4E4E4C4A", x"47464443", x"42424140", x"413F3F41", x"413D3C3D", x"39383A39", x"3B393134",
									 -- x"37363737", x"37353639", x"37353435", x"37383736", x"353A3838", x"3C3A373A", x"3B3C3C3A", x"3B3E4040",
									 -- x"40444545", x"46494A47", x"4B4C5054", x"55535355", x"5858595B", x"5F616160", x"5E646A6A", x"6A6C7173",
									 -- x"76777879", x"7A7B7A79", x"7E7E8081", x"81818284", x"84848380", x"80818281", x"86848385", x"87898888",
									 -- x"8C898B8C", x"8A8C8E8C", x"8E8E8D8C", x"8C8D9092", x"92929191", x"92939495", x"8F939493", x"94989896",
									 -- x"93959798", x"97959494", x"93919092", x"928F8D8C", x"8F8C8987", x"84828182", x"7F7D7D7D", x"79726E6F",
									 -- x"4846494A", x"48484743", x"47444245", x"4B4E4B48", x"4A4B4948", x"47474440", x"403E3C3C", x"3D3D3B38",
									 -- x"3E3D3C3A", x"3837393B", x"35353535", x"36373838", x"33323232", x"322F2D2B", x"2929292A", x"2D323332",
									 -- x"32343636", x"34333436", x"35313034", x"38383635", x"37393A3B", x"3F434543", x"4B4F5355", x"575C5F5F",
									 -- x"60646A6D", x"6F73787C", x"84898E90", x"94999E9F", x"A3A7ABAD", x"ACABAAAB", x"AFAFB0B2", x"B4B7B9BA",
									 -- x"BDC0C1C4", x"C6C3C1C5", x"C2C1C0BF", x"C0C2C3C3", x"C3C4C3C3", x"C4C5C6C6", x"C9C6C6CA", x"CDCED0D3",
									 -- x"D5D5D6D8", x"DDE2E1DC", x"D9DAD9D7", x"D4D3D2D3", x"D0D2D5D9", x"DADCE1E7", x"E5E7E8E7", x"E8EBEEF0",
									 -- x"EFEEECEB", x"ECEFF4F8", x"FAFDFFFE", x"FFFFFFFC", x"EFEAE5E3", x"E3E0DDDB", x"DCE1E1E0", x"E3E1DDDC",
									 -- x"E1E0DDDA", x"D8D8DADC", x"DBDCDFE1", x"E3E5E8E9", x"EEEBE9E8", x"E6E0DAD7", x"D4D3D2D2", x"D4D6D8DA",
									 -- x"DBDAD8D7", x"D7D8DADB", x"DBD8DADD", x"DDE0E2E0", x"E5EBF0F3", x"F7FBF9F3", x"F0EAE9ED", x"ECEAE5DE",
									 -- x"E4E5E7E8", x"E6E4E7EB", x"E8E9E9EA", x"E9E9E8E7", x"E4E5E3DE", x"DBDCDEDE", x"E0E2E4E5", x"E3E1E0E1",
									 -- x"E2E1E0E0", x"E0DEDBD9", x"DEDCDAD7", x"D7D8D5D0", x"D0D3D6D6", x"D4CFCAC7", x"C3C3BEB7", x"B3B3AFAA",
									 -- x"A9A6A4A3", x"A09C9B9C", x"9394928F", x"8D8E8E8E", x"93959799", x"9A9A9B9C", x"9E9E9D9D", x"9C9A9998",
									 -- x"99999993", x"8E939590", x"8F8F8E8D", x"8B898988", x"8A8B8D8E", x"8D898582", x"86858682", x"7F818078",
									 -- x"7D7B7876", x"7573706D", x"6C696967", x"61606364", x"5F605F5F", x"5F5A5657", x"58535053", x"57575351",
									 -- x"534E4C4E", x"4E4B494A", x"46444240", x"3F3E3D3C", x"3D3E3E3D", x"3C3C3B38", x"3B363534", x"393A3234",
									 -- x"37363536", x"35343435", x"34323133", x"35373534", x"35393636", x"3E3D373A", x"3A3B3B3A", x"3C404242",
									 -- x"40424241", x"43484946", x"46484E54", x"54505156", x"59595A5B", x"5C5E5F5F", x"62656768", x"6B6F706E",
									 -- x"74757778", x"7A797876", x"73767C83", x"84818185", x"807F7E7D", x"7F82817E", x"837E7D83", x"86838284",
									 -- x"89868687", x"86888A87", x"8D8C8D8D", x"8E8E8D8C", x"92918F8E", x"8E8F9192", x"8D919291", x"91959694",
									 -- x"94949492", x"908F9192", x"8F8C8B8D", x"8D8B8988", x"88868585", x"827E7B7B", x"78797B7B", x"756C696A",
									 -- x"4B454448", x"49444244", x"45444243", x"46484746", x"43464847", x"423E3C3C", x"3C3B3B3A", x"3A393838",
									 -- x"393B3B38", x"37383939", x"3A393737", x"36353434", x"32343433", x"32312F2C", x"2E2E2D2D", x"2D2E2F30",
									 -- x"30333431", x"30313131", x"32303134", x"35353639", x"36383A3A", x"3C414446", x"4B4E5254", x"575B5E60",
									 -- x"6664656C", x"72757A7F", x"8285898E", x"92979DA0", x"A2A6ACB1", x"B2B0B0B2", x"B2B3B4B4", x"B5B9BBBB",
									 -- x"C0C0C1C2", x"C4C6C7C8", x"C3C1C2C5", x"C8C7C7C8", x"C5C6C6C5", x"C6C9CAC9", x"C7C7C9CC", x"CECFD2D6",
									 -- x"D8D9D9DA", x"DEE1E1DF", x"DDDBDADA", x"DBDBD9D7", x"D6D7D8DB", x"DEE1E4E5", x"E5E6E8E8", x"E8E9EDF0",
									 -- x"F1F2F1EF", x"EEF1F8FE", x"FEFEFEFE", x"FFFEFEFD", x"F0E9E4E3", x"E4E2DFDD", x"D9DDE2E6", x"E6E5E3E2",
									 -- x"E3E2E0DE", x"DFE0E3E5", x"E5E3E2E2", x"E2E3E7EA", x"EAEAEAE8", x"E5E0DCD9", x"D6D4D3D5", x"D6D7D9DB",
									 -- x"DDD9D4D4", x"D6DADBDB", x"DEDBD9DB", x"DCDDDFE2", x"E6E7EAEF", x"F3F5F4F3", x"EFEFEFEE", x"EBE8E4E1",
									 -- x"E4E9EBE7", x"E3E2E5E7", x"EBEAEBEB", x"ECEAE8E5", x"E3E8E7E3", x"E1DEE0E7", x"E4E4E4E5", x"E5E4E2E1",
									 -- x"E2E1E0DF", x"DEDBD7D4", x"D8DADAD8", x"D5D4D4D2", x"CDCECECE", x"CFCFCBC5", x"C0C0BDB8", x"B2ADACAC",
									 -- x"A9A6A6A3", x"9D9B9B98", x"96959391", x"91908C87", x"92929394", x"97999C9D", x"9F9E9C9B", x"99999999",
									 -- x"9A969393", x"918E8F92", x"8E8D8B89", x"8A8B8D8F", x"8C8A8887", x"87878583", x"84828282", x"7F7C7B7C",
									 -- x"79767575", x"726D6C6E", x"65676661", x"5F5F5F5C", x"605D5B5B", x"5A565454", x"52515151", x"504F4F51",
									 -- x"4D4D4C4C", x"4A484543", x"423F3D3C", x"3A393B3F", x"3A3A3A39", x"37363636", x"36353433", x"33343333",
									 -- x"312F3031", x"2F303331", x"36323031", x"32313132", x"33363737", x"37383837", x"36373737", x"3B3F403F",
									 -- x"3E414241", x"42464848", x"464A4E50", x"52555554", x"55555A60", x"605B5A5D", x"60626567", x"686B6D70",
									 -- x"706E6E71", x"75777573", x"7478787C", x"7C797C79", x"7F7C7B7C", x"7B78787A", x"7A7F807C", x"7A7F817F",
									 -- x"83858583", x"84868786", x"858C8E89", x"878B8D8C", x"938D8A8B", x"8F908E8C", x"8C8B8B8E", x"91939392",
									 -- x"94929190", x"908F8E8E", x"8C85878C", x"8A8A8A86", x"85848484", x"817C7979", x"79777777", x"736B6869",
									 -- x"48454447", x"47444243", x"43434343", x"44444240", x"40424443", x"403D3C3C", x"3D3B3836", x"36373737",
									 -- x"383A3A37", x"35353534", x"36363636", x"36363535", x"32343433", x"3333322F", x"302F2E2D", x"2D2E2E2F",
									 -- x"2D2F302F", x"2F313231", x"32313134", x"35343638", x"36383A3B", x"3F45494B", x"4A4E5256", x"585B5E5F",
									 -- x"6766676B", x"70757A7F", x"81858A8E", x"91969BA0", x"AAABAEB2", x"B3B2B2B3", x"B5B7B7B6", x"B7B9BBBB",
									 -- x"BEC0C2C4", x"C7C8C9C9", x"C9C7C7C9", x"CAC9C9C9", x"CBCECECC", x"CACACCCC", x"CDCBCCCF", x"D2D3D4D6",
									 -- x"D9DADBDC", x"DFE2E1DE", x"E0DEDCDB", x"DCDDDEDE", x"DCDDDFE1", x"E5E8EBEC", x"EDEEEEED", x"ECECEEF0",
									 -- x"F3F3F2F1", x"F1F4F9FC", x"FEFEFEFE", x"FFFEFEFD", x"F3ECE6E4", x"E5E4E2E1", x"DCDFE4E8", x"EAE8E5E2",
									 -- x"E4E2DFDE", x"DFE1E4E6", x"E7E6E6E8", x"E8E7E9EB", x"EBEAEAE8", x"E4E0DDDA", x"DFDDDBDB", x"DAD9D9DB",
									 -- x"DBD9D8D8", x"DADDDDDD", x"DEDCDBDC", x"DDDDDEE1", x"E6E7EAED", x"F1F2F1F0", x"EFEEEDEB", x"E8E5E3E2",
									 -- x"E1E5E6E4", x"E1E2E5E6", x"E9E8E8E9", x"EAEAE9E8", x"E7EBE9E5", x"E3E0E0E5", x"E4E4E4E4", x"E4E3E1DF",
									 -- x"E1E0DFDD", x"DAD8D5D3", x"D4D6D8D6", x"D4D2D0CE", x"C9CBCBCB", x"CBCBC8C4", x"C3C1BDB7", x"B1AEADAD",
									 -- x"A6A3A2A1", x"9C9A9A96", x"94928F8E", x"8E8D8C8A", x"90909092", x"94979B9D", x"9E9D9C9A", x"98969594",
									 -- x"97949190", x"908E8E8F", x"8C8C8C8C", x"8D8D8D8D", x"8A878584", x"8483807E", x"83818080", x"7E7A7879",
									 -- x"75737272", x"6F6C6B6B", x"63666560", x"5D5E5E5C", x"5B585657", x"56535252", x"504F4E4E", x"4D4C4D4E",
									 -- x"4A494746", x"44423F3D", x"3E3C3B3A", x"3937383A", x"36353433", x"32313131", x"302F2F2F", x"30303030",
									 -- x"31303334", x"3030312F", x"32302F31", x"31323438", x"35363635", x"36383836", x"36363535", x"383C3E3D",
									 -- x"3A3D3F40", x"42454848", x"46494B4B", x"4B4E504F", x"55565757", x"595C5E5E", x"5B5D5F61", x"63666A6D",
									 -- x"6A6A6B6D", x"6E707171", x"6E727175", x"76747977", x"7B787778", x"79787878", x"74767777", x"77797C7E",
									 -- x"81817F7C", x"7D808384", x"858B8D8A", x"8A8D8C87", x"8E8B8A8C", x"8C8B8B8C", x"8E8D8D8D", x"8E8E8C8A",
									 -- x"8F8E8C8B", x"8B8A8988", x"8D888888", x"85838484", x"837F7C7A", x"78767677", x"75727171", x"706C6866",
									 -- x"45454544", x"44434242", x"3F404142", x"413F3D3B", x"3E3E3F3E", x"3C3B3A3A", x"3B393634", x"34343535",
									 -- x"33353634", x"34343433", x"33343636", x"37363535", x"33343433", x"33333331", x"3231302F", x"2E2D2D2D",
									 -- x"2B2B2C2C", x"2E313231", x"33323234", x"34343537", x"383A3C3E", x"41484D4F", x"4B4E5358", x"5A5C5D5F",
									 -- x"67696A6B", x"6E757B7E", x"8185898D", x"90949A9F", x"A8A8AAAF", x"B3B5B7B9", x"B9BBBBB9", x"B9BBBBBB",
									 -- x"BEC0C4C7", x"CACCCDCD", x"D0CECECE", x"CFCDCCCD", x"CED2D2CF", x"CBCACCCD", x"D1CFCFD2", x"D6D7D7D8",
									 -- x"DADCDEE0", x"E3E5E3E0", x"E4E4E3E1", x"E1E1E3E5", x"E2E3E5E7", x"EAEDF0F1", x"F5F5F5F4", x"F1F0F0F0",
									 -- x"F6F5F5F5", x"F7F9FBFC", x"FEFEFEFE", x"FFFEFEFD", x"F5EEE6E3", x"E3E3E2E1", x"E1E2E5E9", x"ECECE9E6",
									 -- x"E6E3E0DF", x"E1E4E6E6", x"E4E5E7EB", x"ECEBEAEA", x"ECECEAE8", x"E5E2DFDE", x"DFDDDDDE", x"DEDDDDDE",
									 -- x"DCDDDEE0", x"E1E1E0E0", x"DFDEDFE0", x"DFDEDEDF", x"E7E8EAEE", x"F2F4F3F2", x"F2F0EDEA", x"E7E6E5E5",
									 -- x"E0E2E3E1", x"E1E2E5E6", x"E7E6E7E8", x"EAEBEAEA", x"EBEDEAE6", x"E5E2E0E3", x"E1E1E2E2", x"E2E1DFDE",
									 -- x"DFDEDDDA", x"D6D3D2D1", x"CDD0D3D2", x"D0CECAC7", x"C5C6C7C7", x"C7C6C5C3", x"C2BEB9B3", x"AFACAAAA",
									 -- x"A4A09F9E", x"9B999893", x"928F8D8D", x"8D8B8C8F", x"94949494", x"94959696", x"95959594", x"94949494",
									 -- x"95949190", x"9192918E", x"8C8C8C8D", x"8D8D8D8D", x"89878583", x"82807D7B", x"7F7D7C7C", x"7B787574",
									 -- x"6F706F6D", x"6B6A6967", x"6164645F", x"5D5D5D5B", x"56545252", x"51505051", x"4E4C4B4A", x"4948494A",
									 -- x"47464442", x"403E3C3B", x"39393839", x"37343334", x"33312F2E", x"2D2D2D2D", x"2D2C2B2B", x"2C2C2D2D",
									 -- x"2F2F3435", x"312F302E", x"2F2F2F2F", x"2F313539", x"37363433", x"35373734", x"35353434", x"363A3B3B",
									 -- x"3B3D3E3E", x"3F424343", x"47494B4A", x"4A4C5051", x"54565452", x"555B5E5B", x"5D5E5E5D", x"5E606467",
									 -- x"67696A69", x"68696C6F", x"6B6E6C6F", x"70707675", x"73737271", x"73757574", x"72717274", x"7575787C",
									 -- x"7A7A7978", x"7A7F8385", x"85858380", x"848C8E8B", x"8B8B8D8C", x"8986888B", x"8B8B8B8C", x"8C8B8A89",
									 -- x"8B8A8988", x"88878685", x"86878482", x"817D7C80", x"7F7C7B7B", x"7A777473", x"73716E6D", x"6E6E6A64",
									 -- x"42444542", x"41424241", x"3B3D3E3E", x"3D3C3B3B", x"3C3C3B3A", x"3A383737", x"35353535", x"34343231",
									 -- x"30323232", x"32343433", x"34363636", x"35353433", x"33343432", x"32333231", x"34333230", x"2F2E2E2E",
									 -- x"2C2B2B2C", x"2F313231", x"34343434", x"34343638", x"3D3F4040", x"43484C4E", x"4D505459", x"5B5C5E60",
									 -- x"656A6D6D", x"6F767B7D", x"8183878B", x"9094999C", x"A2A4A7AD", x"B2B5BABE", x"BCBEBFBD", x"BCBCBDBC",
									 -- x"C1C2C5C8", x"CCCFD1D2", x"D3D2D2D2", x"D2D2D2D2", x"CFD2D3D0", x"CDCDCECF", x"D2D1D2D5", x"D8D8DADB",
									 -- x"DEE0E3E5", x"E8EAEAE7", x"E9EBECEB", x"E9E8E8E9", x"E9EAEBED", x"EFF1F3F3", x"F7F7F8F7", x"F5F3F3F3",
									 -- x"F8F8F9FA", x"FBFCFCFD", x"FEFEFEFE", x"FFFEFEFD", x"F7F0E8E2", x"E1E0DFDE", x"E4E5E6E9", x"EBECEBEB",
									 -- x"E6E4E3E3", x"E6E7E7E7", x"E0E1E6EB", x"EEEDECEC", x"EEEDEBE9", x"E6E5E3E3", x"DDDDDFE3", x"E4E3E3E4",
									 -- x"DFE1E4E6", x"E5E3E1E1", x"E1E2E3E4", x"E2E1E0E0", x"E4E6E9EE", x"F4F6F7F6", x"F4F2EEEB", x"E9E8E8E8",
									 -- x"E2E2E1E0", x"E0E2E4E4", x"E6E7E8EA", x"EBEBEBEA", x"EBEBE8E5", x"E5E2DFE1", x"DFDFDFE0", x"E0DFDDDC",
									 -- x"DADAD9D7", x"D3D0CECE", x"C7CACCCC", x"CAC8C5C1", x"C1C3C4C3", x"C2C2C2C2", x"C0BCB6B1", x"AEACA9A7",
									 -- x"A39F9E9E", x"9B999792", x"938E8C8E", x"8D8A8C92", x"94949595", x"94939190", x"908F8F8F", x"91939698",
									 -- x"93939290", x"9194928D", x"8E8D8B89", x"89898B8C", x"88868483", x"817F7C7A", x"7A787777", x"78767370",
									 -- x"6C6E6D69", x"68686662", x"6062615F", x"5E5F5C58", x"5452504F", x"4F4F4F4F", x"4E4B4847", x"46454546",
									 -- x"4342403F", x"3E3E3D3C", x"38373737", x"35323030", x"31302E2D", x"2D2D2D2C", x"2E2C2A2A", x"2A2B2C2D",
									 -- x"2C2D3234", x"2F2F302F", x"2F2F2F2F", x"2F303235", x"35353432", x"32343432", x"32343434", x"36383A39",
									 -- x"3A3B3D3D", x"3E3F4041", x"47494B4B", x"4B4E5255", x"52545553", x"55585958", x"5F5E5D5B", x"5B5D6165",
									 -- x"66676867", x"6565686A", x"696C696C", x"6D6C7271", x"6D70706D", x"6D70716F", x"71717172", x"72737679",
									 -- x"74757678", x"7B7E8081", x"81807B79", x"7D868A89", x"8B8C8E8C", x"8884868B", x"8788898A", x"8A898988",
									 -- x"86878786", x"86878583", x"7C807D7B", x"7E7B787C", x"76757677", x"75716E6D", x"72716D6A", x"6A6C6862",
									 -- x"40434440", x"3F424340", x"3C3C3B3A", x"393A3B3D", x"3A3A3A39", x"38363433", x"32323233", x"33333230",
									 -- x"33333230", x"2F313231", x"33353533", x"32333332", x"33343432", x"32343433", x"34343332", x"32313130",
									 -- x"2F2D2D2F", x"31333434", x"35363736", x"3637393B", x"41424342", x"44484B4D", x"5152565A", x"5C5D5F63",
									 -- x"636A6E6F", x"72777B7C", x"8182858A", x"9096999A", x"A1A5AAAE", x"B0B3B8BE", x"BDC0C1C0", x"BEBEBFBE",
									 -- x"C3C4C5C7", x"CBCFD3D5", x"D3D3D4D4", x"D5D6D6D6", x"D3D5D5D4", x"D3D4D4D3", x"D4D5D8DA", x"DADADCDF",
									 -- x"E4E7E9EA", x"EDEFEFEE", x"EEF0F2F1", x"EFEEEFF0", x"F3F3F4F5", x"F6F6F7F7", x"F5F6F8F8", x"F8F8F8F8",
									 -- x"FAFBFDFE", x"FDFCFDFE", x"FEFEFEFE", x"FFFEFEFD", x"F8F3EBE5", x"E2E1E0DE", x"E4E7EAEB", x"EAE8E8E9",
									 -- x"E4E5E6E8", x"E9EAE8E7", x"E1E2E5EA", x"EEEEEEEE", x"EDECEAE9", x"E7E7E6E6", x"E4E4E8EB", x"EDEBE9E9",
									 -- x"E5E7EAEA", x"E8E5E3E3", x"E4E6E7E7", x"E6E4E3E1", x"E0E2E6EC", x"F2F6F6F6", x"F3F1EFED", x"EBEAE9E9",
									 -- x"E6E3E1E0", x"E0E1E1E1", x"E6E7EAEB", x"ECEBE9E8", x"E7E8E4E2", x"E4E3E0E1", x"DFDFDFDF", x"DEDDDBD9",
									 -- x"D4D5D5D3", x"D0CDCBC9", x"C6C7C8C7", x"C6C5C2BF", x"C0C0C0C0", x"BFBFC0C1", x"BEBBB6B3", x"B1AEAAA7",
									 -- x"A39F9E9E", x"9C9B9994", x"928E8C8E", x"8D898B90", x"8E8E8F8F", x"8F8F8E8E", x"90909090", x"91929293",
									 -- x"9091908E", x"90928F8A", x"8C8B8886", x"85858586", x"84838180", x"7E7D7B7A", x"79777574", x"7473706D",
									 -- x"6A6C6A66", x"6566635F", x"5D5E5D5C", x"5D5E5952", x"5352504E", x"4E4D4D4C", x"4D494645", x"43424142",
									 -- x"3F3D3C3B", x"3B3B3B3A", x"38363535", x"33302E2E", x"2F2F2E2E", x"2E2D2B2A", x"2F2D2A29", x"2A2C2E30",
									 -- x"2C2D3132", x"2F2F3130", x"30303030", x"31323130", x"31333432", x"2F2F3030", x"30333535", x"37383938",
									 -- x"3637393C", x"3E404244", x"45474849", x"494A4D50", x"4F505356", x"54525458", x"58585757", x"585B6063",
									 -- x"61626363", x"63636464", x"65686568", x"6A696D6C", x"6A6E706C", x"6A6C6D6D", x"6B6E6F6C", x"6D727473",
									 -- x"74747577", x"78797B7C", x"7C7E7E7D", x"7E80807E", x"8A898988", x"8685868A", x"87888887", x"85838282",
									 -- x"81838382", x"8182807D", x"7B7D7775", x"7A797678", x"76747371", x"6E6C6D70", x"6A6B6964", x"6364625E",
									 -- x"41424240", x"40424341", x"3F3D3A38", x"37383A3B", x"38393938", x"35333231", x"32312F2F", x"30313232",
									 -- x"32312F2D", x"2E313231", x"2E32322F", x"2F313332", x"33343434", x"34373737", x"35343434", x"34333333",
									 -- x"32303033", x"3536383A", x"37393A39", x"383B3E40", x"43454545", x"464A4D4D", x"5454575C", x"5E5E6165",
									 -- x"65696E71", x"74787B7C", x"8183868C", x"91969899", x"9EA2A9AD", x"AEB0B6BD", x"BFC2C4C3", x"C1C1C1C1",
									 -- x"C4C5C6C8", x"CBCED2D4", x"D2D5D6D7", x"D7D8D8D8", x"D8D9D9D8", x"D9DADAD8", x"DADCDFE0", x"DEDDDFE3",
									 -- x"EBEDEFEF", x"F0F2F2F0", x"F2F2F3F2", x"F1F3F6F9", x"F9F9F9FA", x"FAFAF9F9", x"F6F7F9FA", x"FCFCFDFD",
									 -- x"FBFDFFFF", x"FEFDFDFF", x"FEFEFEFE", x"FFFEFEFD", x"F7F3EDE7", x"E5E4E1DF", x"E2E7EDEE", x"EAE6E3E3",
									 -- x"E3E4E6E7", x"E8E8E8E7", x"E5E3E4E7", x"EAEAEAEB", x"EAEAEAE9", x"E9E8E8E8", x"E8E9ECEF", x"F1EFEEEE",
									 -- x"EDEFF1F1", x"EEEBE9E8", x"E8E9E9E8", x"E8E7E4E1", x"E0E2E5EB", x"F0F3F3F2", x"F2F1F0EF", x"EDECECEB",
									 -- x"EAE7E4E3", x"E2E1E0E0", x"E3E5E9EA", x"EAE8E6E5", x"E3E4E0DF", x"E2E1DFE0", x"E0E0DFDE", x"DCD9D6D4",
									 -- x"D0CFCFCE", x"CDCAC7C4", x"C4C5C4C2", x"C1C1C0BE", x"BEBCBBBB", x"BBBBBCBE", x"B9B7B4B2", x"B0AEAAA6",
									 -- x"A29E9F9F", x"9D9C9C98", x"918D8B8B", x"8A88888B", x"8F8E8B89", x"89898B8C", x"888A8C8E", x"8F8E8C8B",
									 -- x"90908F8E", x"8F8F8D89", x"87878685", x"83817F7E", x"81807F7D", x"7C7B7A7A", x"79787673", x"71706D6A",
									 -- x"69686663", x"62625F5D", x"595A5857", x"595A544C", x"50504F4D", x"4C4B4946", x"49464242", x"413F3E3E",
									 -- x"3D3C3A39", x"39383837", x"37353333", x"322F2D2D", x"2B2C2D2D", x"2C2A2929", x"2D2B2A29", x"2B2D2F31",
									 -- x"2F2D3031", x"2F303230", x"31313131", x"33353330", x"2E323431", x"2D2D2E2F", x"2F323435", x"36373737",
									 -- x"3737393B", x"3D3F4144", x"46454647", x"46454547", x"4C4C4F53", x"514E5259", x"55555656", x"56585B5E",
									 -- x"5C5C5E60", x"62636261", x"62646266", x"69686C6A", x"686C6E6D", x"6A6A6B6B", x"676C6D69", x"6B727470",
									 -- x"74737375", x"77797C7E", x"7A7D7E7C", x"7C7E7F7F", x"83818182", x"83848586", x"82848482", x"7F7D7D7E",
									 -- x"7F81817E", x"7D7D7975", x"7F7D7671", x"74757474", x"74737272", x"6F6C6C6D", x"63656462", x"5F5F5F5E",
									 -- x"42414040", x"41434342", x"403D3A38", x"38393938", x"36373735", x"32313233", x"302F2E2E", x"2F2F3030",
									 -- x"2E2E2D2B", x"2D303130", x"2C30322F", x"2F313332", x"32343534", x"35383838", x"34343535", x"34343434",
									 -- x"36353537", x"3737393D", x"393C3D3C", x"3B3F4345", x"45474848", x"4A4D4F4F", x"5656595E", x"605F6166",
									 -- x"68696D72", x"76787A7B", x"82868B90", x"92959799", x"9C9FA5AA", x"ADB0B7BE", x"C0C5C7C6", x"C4C3C3C3",
									 -- x"C5C7C9CD", x"CFD0D1D1", x"D1D5D8D9", x"D9DBDCDB", x"D9DBDDDC", x"DCDEDEDE", x"E0E1E3E5", x"E4E2E4E7",
									 -- x"ECEFF2F2", x"F3F4F3F1", x"F2F3F3F3", x"F3F5F9FB", x"F9FAFBFB", x"FCFCFBFB", x"FAFAFAFC", x"FDFEFEFE",
									 -- x"FEFEFEFE", x"FEFEFEFD", x"FEFEFEFE", x"FFFEFEFD", x"F8F6F2ED", x"EAE8E4DF", x"E2E6EAEC", x"E9E5E3E2",
									 -- x"E2E3E3E3", x"E2E3E6E9", x"E8E5E3E5", x"E7E7E7E8", x"E9E9EAEB", x"EBEBEBEB", x"E8E8E9EC", x"EDEDEEF0",
									 -- x"EFF1F3F4", x"F3F0EEEC", x"EAEAE8E6", x"E7E7E4DF", x"E0E1E4E8", x"ECEEEEEC", x"EEEEEDEC", x"ECEBEBEB",
									 -- x"EAE7E4E4", x"E2E0DEDF", x"DEE1E4E5", x"E5E3E2E2", x"DEDFDBD9", x"DCDCDADC", x"DCDCDBD9", x"D7D5D1CF",
									 -- x"CDCBC9C8", x"C8C6C2BF", x"C1C0BEBC", x"BCBDBCBA", x"BBB7B4B5", x"B6B6B7B9", x"B4B2B1B0", x"AEACA9A6",
									 -- x"A2A0A0A0", x"9C9B9B98", x"918E8A88", x"87878787", x"8F8D8A87", x"86868687", x"82848689", x"8A8B8A8A",
									 -- x"908F8E8F", x"8E8C8989", x"84848382", x"807E7C7A", x"7D7D7B79", x"78787879", x"7576736F", x"6D6D6B69",
									 -- x"6763605F", x"5F5D5C5B", x"57585653", x"5354514C", x"4D4E4E4C", x"4B4A4642", x"44413E3E", x"3F3D3C3C",
									 -- x"3D3C3A39", x"38373635", x"33313031", x"312F2D2C", x"2A2D2E2D", x"2B29292A", x"2C2B2B2B", x"2C2D2E2E",
									 -- x"2D2B2D2F", x"2E30312E", x"2F313231", x"32343331", x"2F31312E", x"2C2C2E2E", x"2F313332", x"32343535",
									 -- x"3A39393B", x"3C3C3F42", x"46434244", x"45444445", x"484A4C4D", x"4C4C4F53", x"54555656", x"55555657",
									 -- x"59595B5D", x"5F605F5E", x"60626064", x"66666967", x"6565676A", x"6A696868", x"67696B6A", x"6D70716F",
									 -- x"72717275", x"77787A7D", x"78797877", x"787C8082", x"7D7B7B7E", x"81818181", x"7D7F807F", x"7C7B7D7F",
									 -- x"7D807F7C", x"7A797570", x"7B787571", x"6F70716E", x"6C6A6A6C", x"6C686361", x"61616262", x"605D5D5F",
									 -- x"44413F40", x"43434342", x"3E3C3A39", x"3A3A3836", x"34353533", x"30303235", x"2D2D2E2F", x"302F2D2C",
									 -- x"2F2E2D2B", x"2C2E2D2B", x"2C323431", x"30333331", x"32343534", x"35363735", x"34343535", x"35343434",
									 -- x"3A39393A", x"3837393D", x"393D3F3D", x"3D414648", x"474A4B4B", x"4C4F5050", x"56565A61", x"62606166",
									 -- x"6B6A6C73", x"7777797C", x"82889093", x"9393979A", x"A1A2A5AA", x"AEB2B8BE", x"C2C6C9C8", x"C5C5C5C5",
									 -- x"C6C9CED2", x"D4D3D1D0", x"D0D5D9DA", x"DBDEDFDE", x"D9DEE1E1", x"E0E1E3E5", x"E2E2E4E7", x"E7E7E7E9",
									 -- x"EBEFF2F4", x"F4F5F3F1", x"F1F2F4F5", x"F6F7F7F8", x"FAFAFCFD", x"FEFEFEFE", x"FCFCFCFC", x"FCFDFCFC",
									 -- x"FFFEFDFD", x"FFFFFEFC", x"FEFEFEFE", x"FFFEFEFD", x"FDFCF8F3", x"EFECE7E1", x"E3E4E5E7", x"E7E6E6E6",
									 -- x"E1E1E0DE", x"DCDFE5EA", x"EBE7E5E6", x"E8E8E8E9", x"E9EAECED", x"EEEEEEEE", x"EBE9E8E8", x"E9E8EAEC",
									 -- x"EBEDF0F2", x"F2F0EDEA", x"ECEAE7E5", x"E6E6E2DD", x"DDDEE0E4", x"E7E9E8E7", x"E8E8E7E6", x"E6E6E6E6",
									 -- x"E5E2E0E0", x"DFDCDADB", x"DADCDFE0", x"E0E0E0E1", x"DADBD7D5", x"D7D7D6D8", x"D6D6D5D4", x"D3D1CECC",
									 -- x"CDC9C5C4", x"C5C3BFBB", x"BCBCBAB8", x"B8B9B8B5", x"B9B4B0B1", x"B2B3B4B5", x"B2B2B1AF", x"AEACAAA9",
									 -- x"A4A1A2A0", x"9A999997", x"928F8A85", x"85888886", x"87878787", x"86848383", x"86868586", x"87898B8C",
									 -- x"8F8C8B8D", x"8B878587", x"8482807E", x"7C7B7B7B", x"79787674", x"73737475", x"7071706C", x"696A6A69",
									 -- x"655F5C5D", x"5D5B595B", x"56585752", x"4F50504E", x"4B4D4E4C", x"4B494540", x"403D3B3C", x"3D3C3A3A",
									 -- x"3A393837", x"37363534", x"302E2E30", x"312F2C2C", x"2C2F302E", x"2B292B2D", x"2D2D2D2D", x"2D2D2B2A",
									 -- x"2927292D", x"2E30312D", x"2E313230", x"2F303231", x"31312F2C", x"2B2D2E2E", x"2F313130", x"2F313334",
									 -- x"3937373A", x"3B3C4044", x"433F3E41", x"44454547", x"43494C4A", x"4A4D4C49", x"4E505354", x"54545555",
									 -- x"55565758", x"59595858", x"5F605C5F", x"61606462", x"625F6066", x"6A686564", x"6867686B", x"6D6C6C6D",
									 -- x"71707276", x"76737172", x"73747677", x"78797978", x"7A797A7D", x"7F7E7D7C", x"7D7F807E", x"7A797C7F",
									 -- x"797C7C78", x"7776726C", x"72717473", x"6D6E7069", x"726B6666", x"69686562", x"615F5F61", x"605C5B5E",
									 -- x"40424240", x"3E3E3E3D", x"383C3E3C", x"38363331", x"33363835", x"2F2C2E32", x"2D2E2C2A", x"2B2D2E2C",
									 -- x"29292A2A", x"2827292D", x"292A2D30", x"32323335", x"32343434", x"34363635", x"36343233", x"34343538",
									 -- x"38393A3B", x"3B3A3A3A", x"3E3D3D3F", x"43464646", x"4B4A4A4B", x"4F525353", x"555C5D5C", x"6060636C",
									 -- x"6868686E", x"7779787B", x"84898B8D", x"9295979D", x"A0A7A9AA", x"B0B1B6C3", x"C7C8C8C7", x"C6C6C8C9",
									 -- x"CACCD0D3", x"D6D6D6D6", x"D3D7DADB", x"DCDFE0E0", x"DFDFE2E7", x"EBEDEAE7", x"E8E4E3E5", x"E8EBECEE",
									 -- x"EDEEF0F0", x"F0F0F0EF", x"F2F5F4F2", x"F4F4F6FB", x"F9FBFEFF", x"FEFDFEFE", x"FCFCFDFD", x"FEFEFEFD",
									 -- x"FFFFFEFE", x"FFFFFFFE", x"FFFFFEFC", x"FAFBFEFF", x"FDFBF6EF", x"EDEEEDEC", x"E9E6E5E6", x"E7E5E5E7",
									 -- x"E2DEDBDB", x"DCDCE2EA", x"E9E9E9EA", x"ECECECEB", x"EAE9EBF0", x"F2F2F2F2", x"EFEAE7E6", x"E6E4E4E6",
									 -- x"E4E6E9EC", x"EDECEBEA", x"EEEBE8E6", x"E6E5E1DB", x"DADDE0E1", x"E2E2E1DF", x"DFE0E0DF", x"DFE1E1E0",
									 -- x"E1DDDBDA", x"D9D7D7D8", x"D7D7D8DA", x"DCDEDBD8", x"DAD5D2D1", x"D1CFCFD0", x"D0CFCFCE", x"CDCBC9C7",
									 -- x"C6C5C2BF", x"BDBAB8B7", x"BBB7B4B3", x"B3B3B0AC", x"B1B3AFAB", x"ACADACAD", x"B3B1AFAD", x"ABAAA9A8",
									 -- x"A4A19E9B", x"99989594", x"938F8A86", x"83828487", x"8482807D", x"7D7D7D7C", x"7C7D7E80", x"8386888A",
									 -- x"89878689", x"89868382", x"7F7D7D7C", x"7A767678", x"77747171", x"72716E6A", x"6868696A", x"6966625F",
									 -- x"615E5B59", x"5A595856", x"5454524F", x"4E4E4D4A", x"4C494848", x"47444343", x"3A3B3B39", x"3A3C3A36",
									 -- x"34353534", x"3434322F", x"2E302F2D", x"2E312E29", x"2C2D2F2F", x"2D2C2B2B", x"2D2C2B2A", x"2B2D2D2C",
									 -- x"292C2D2B", x"2C2E2F2C", x"2D2E2E2C", x"2C2D2D2B", x"342F2B2A", x"2E302F2C", x"2A2F2D2A", x"2F353635",
									 -- x"3A383537", x"3B3A3A40", x"40404345", x"44424245", x"4A484747", x"48494A4A", x"4C4F5151", x"4E4D5052",
									 -- x"50545859", x"57555557", x"5B5B5A5A", x"5B5D5F61", x"5F63615E", x"62646261", x"696A6864", x"656B6F6F",
									 -- x"6B6E7071", x"71737372", x"71737576", x"76777572", x"7B77767A", x"7B78797E", x"7A7A7B7C", x"7A767779",
									 -- x"75737577", x"7371706D", x"6D71726E", x"6A696B6C", x"6A686462", x"61616263", x"5F635F5B", x"5D5B595F",
									 -- x"3D40403E", x"3C3C3D3C", x"3A3C3C3A", x"37373634", x"32323231", x"2F2D2D2E", x"292B2C2C", x"2D2E2D2A",
									 -- x"27272728", x"2726292D", x"2A292B2E", x"30303133", x"32343332", x"33353636", x"37353536", x"3636383B",
									 -- x"3A3B3D3D", x"3C3B3B3B", x"3E3D3C3D", x"40434545", x"4B4B4C4E", x"50525556", x"575A5B5D", x"6264666A",
									 -- x"6B6C6C70", x"787A7A7E", x"81878B8E", x"9395979C", x"A2A9AAAD", x"B2B3B7C1", x"C7C9CAC9", x"C7C7C9CB",
									 -- x"D0D1D2D4", x"D5D6D7D7", x"DBDCDDDE", x"E0E3E3E1", x"E2E3E5E9", x"EDEEECEA", x"E9E6E6E9", x"ECEDEEEF",
									 -- x"F0F0EFEE", x"EDECEBEB", x"EDF0F0EF", x"F2F2F4F9", x"F9F9FAFB", x"FCFDFCFC", x"FDFDFDFD", x"FDFEFFFF",
									 -- x"FFFFFFFF", x"FFFFFEFD", x"FFFDFAF9", x"FAFBFCFC", x"FBFBF9F4", x"F2F2F1EF", x"EEEBEAEB", x"EAE7E5E5",
									 -- x"DFDAD7D7", x"D7D8DFE6", x"E7E8E9EC", x"EEF0EFEE", x"EDEBEBEF", x"F3F4F2F2", x"ECEAE8E9", x"E8E5E2E1",
									 -- x"E5E6E6E6", x"E7E8E9E9", x"EBEBE9E6", x"E5E4E2DE", x"DBDDDDDC", x"DCDDDDDB", x"DADBDBD9", x"D9DBDBDA",
									 -- x"DDDAD9D9", x"D8D6D4D5", x"D1D1D2D4", x"D6D6D4D2", x"D4D0CDCD", x"CECDCDCE", x"CDCCCBCA", x"C9C6C4C2",
									 -- x"BFBDBAB9", x"B8B6B5B3", x"B5B2B0AF", x"B0B0ADAB", x"ABAFADA9", x"AAAAAAAD", x"ACABAAA9", x"A7A6A5A5",
									 -- x"A4A19E9B", x"99969391", x"8F8B8684", x"83838485", x"8381807E", x"7E7D7B7A", x"797A7B7D", x"80828485",
									 -- x"89868484", x"84817E7E", x"7C7B7A7A", x"78747476", x"71706E6D", x"6E6D6A68", x"68676562", x"5E5B5A5A",
									 -- x"5B585553", x"5353514F", x"4F4F4D4B", x"4A494845", x"45434241", x"403D3C3D", x"3A3A3937", x"37383735",
									 -- x"36343231", x"302F2E2D", x"2D2D2D2D", x"2E2F2D2A", x"2B2D2E2E", x"2D2C2D2E", x"2F2E2E2E", x"2E2C2B2A",
									 -- x"292B2C2B", x"2B2C2E2E", x"2D2D2B2A", x"2C2E2C29", x"312E2C2C", x"2F302F2D", x"292E2D2C", x"31353535",
									 -- x"35363537", x"3C3C3B3F", x"3E3E3F43", x"44434243", x"43434546", x"47484848", x"4A4C4E50", x"50505051",
									 -- x"4F525556", x"56555556", x"57575657", x"585A5B5D", x"5E605E5D", x"61636263", x"65676764", x"656A6D6B",
									 -- x"6E70706F", x"6E6D6D6B", x"71747675", x"74747372", x"78787776", x"77797A7A", x"7A79797A", x"79767575",
									 -- x"74727373", x"706F6F6C", x"6A6D6D69", x"66666767", x"68666362", x"615F5C5A", x"5E61605E", x"5C585556",
									 -- x"3E3F3F3C", x"3A3B3B3B", x"393A3A39", x"39383734", x"312F2C2C", x"2E2F2D2A", x"2A2B2C2C", x"2D2D2C2A",
									 -- x"27262626", x"2625282C", x"2C29292B", x"2D2D2E2F", x"31323231", x"32363838", x"38373738", x"38383A3E",
									 -- x"3A3D3F3F", x"3E3D3D3E", x"40404040", x"4144484A", x"4B4D5051", x"51535659", x"5A585B5F", x"63676A68",
									 -- x"6D6F6E71", x"77787A7F", x"80868B8F", x"9496989D", x"A2A7AAAE", x"B4B5B8BF", x"C6C8CBCB", x"C9C9CDD0",
									 -- x"D3D4D4D4", x"D4D5D7D8", x"DFDEDDDE", x"E1E4E3DF", x"E3E5E7E9", x"EBECECEC", x"E9E8E9ED", x"F0F1F1F2",
									 -- x"F3F2F1EE", x"ECEAE9E8", x"E8EBEBEB", x"EFF1F2F7", x"F9F8F8FA", x"FCFEFDFB", x"FCFCFCFC", x"FCFEFFFF",
									 -- x"FFFFFFFF", x"FFFEFDFC", x"FEFAF7F8", x"FCFEFCFA", x"F7F9FAF7", x"F5F3F2F1", x"F1EFEDEE", x"EDEAE6E3",
									 -- x"DDD9D5D4", x"D4D6DBE1", x"E3E5E8EB", x"EFF1F1F1", x"EFEBEAED", x"F2F3F1EF", x"EDEBEAEB", x"EAE6E2E0",
									 -- x"E5E4E4E3", x"E4E5E6E7", x"E9EAE9E5", x"E3E2E2E0", x"DDDDDBD8", x"D7D8D8D7", x"D5D7D7D5", x"D5D6D6D5",
									 -- x"D5D4D3D4", x"D4D1CFCE", x"CECCCDD0", x"D2CFCDCE", x"CECBC8C8", x"C8C8C8C8", x"C9C8C6C4", x"C2C0BDBB",
									 -- x"B9B7B4B3", x"B3B3B1AF", x"AFAEACAC", x"ACABAAA9", x"A4A9A8A5", x"A5A5A5A9", x"A4A4A3A3", x"A2A1A1A0",
									 -- x"9F9D9B99", x"9794918E", x"8A868282", x"83838281", x"7F7E7E7E", x"7D7B7877", x"77787A7C", x"7F808182",
									 -- x"86827F7E", x"7D7B7A79", x"79787877", x"74716F70", x"6D6C6B6A", x"69676564", x"62615F5B", x"58565759",
									 -- x"55524F4E", x"4D4D4C4A", x"4A4A4947", x"47464442", x"413F3E3D", x"3B383839", x"38383735", x"33343434",
									 -- x"35312E2E", x"2E2B2C2E", x"2E2C2C2F", x"302F2E2D", x"2A2C2E2E", x"2C2C2E30", x"2C2C2E31", x"302C2A2B",
									 -- x"2B2B2B2B", x"2A2A2C2F", x"2F2D2B2B", x"2F312F2A", x"2F2F2F30", x"3131302E", x"2A2D2D2F", x"33343234",
									 -- x"32363738", x"3C3D3B3B", x"3A393B3F", x"42424141", x"40414445", x"45464748", x"48494B4E", x"4F4F4E4D",
									 -- x"4E4F5152", x"53545453", x"54545556", x"57585A5A", x"5B5C5A5B", x"5F605F63", x"61646565", x"66696967",
									 -- x"696C6D6C", x"6C6D6D6C", x"70747573", x"70717273", x"74797871", x"71777974", x"76747374", x"7472706F",
									 -- x"706D6E6D", x"6A6B6C6A", x"67686765", x"63636261", x"6362605F", x"5E5B5855", x"5D5C5E5E", x"59555350",
									 -- x"4041403D", x"3A3A3B3B", x"39393B3D", x"3E3C3833", x"332F2B2B", x"2E2F2C28", x"2E2D2B2A", x"2A2B2B2A",
									 -- x"29272626", x"25252629", x"2C292729", x"2B2B2B2B", x"2F313131", x"33373A3A", x"37383939", x"38383B3D",
									 -- x"3A3D4041", x"403F3F41", x"3F414243", x"44464B4E", x"4E4F5152", x"53555759", x"5C595D61", x"61686D68",
									 -- x"6E707173", x"7778797F", x"81888C8F", x"95979A9F", x"A1A4A9AF", x"B5B7B9BD", x"C2C7CBCC", x"CACBD0D4",
									 -- x"D3D5D6D6", x"D6D7D8D9", x"DEDEDDDD", x"DFE1E1DF", x"E2E3E6E7", x"E7E7E8E9", x"E8E7E9ED", x"F1F3F4F5",
									 -- x"F4F3F1F0", x"EDEBE9E7", x"E3E6E5E6", x"EBEEEEF2", x"F6F6F6F8", x"FAFCFCFC", x"FAFAFAFB", x"FCFDFEFF",
									 -- x"FEFEFFFF", x"FFFEFCFA", x"FAF8F6F8", x"FCFDFBF8", x"F5F7F8F7", x"F4F2F2F2", x"F2F0EEEE", x"EEEBE7E4",
									 -- x"DFDBD8D7", x"D7D7DADE", x"E0E2E5E8", x"EBEEEFEF", x"EDEBEAEB", x"EEF0EEED", x"EDECEAE9", x"E9E7E4E2",
									 -- x"E2E3E4E5", x"E6E5E5E4", x"E8E9E7E3", x"E1E1E0DF", x"DFDFDCD8", x"D6D5D5D4", x"D2D4D4D3", x"D2D3D3D2",
									 -- x"D0CFCFD0", x"CFCECCCB", x"CCC9C9CD", x"CECBCACB", x"CAC7C4C3", x"C3C3C2C2", x"C4C2C1BF", x"BDBBB8B7",
									 -- x"B5B2AFAE", x"AFAEABA9", x"A9A9A8A7", x"A6A4A4A3", x"A0A3A2A0", x"A1A09FA1", x"9F9F9F9F", x"9F9E9D9C",
									 -- x"98979695", x"94918E8B", x"88848282", x"82807E7D", x"7C7B7A7B", x"79767474", x"76787A7C", x"7E7F7F7F",
									 -- x"7F7D7B7A", x"79787777", x"77767573", x"706D6A6A", x"69686765", x"62605E5D", x"59595958", x"56555555",
									 -- x"504E4C4B", x"4B4B4A4A", x"44454544", x"4343423F", x"3F3D3B3B", x"3A383635", x"35363634", x"32313233",
									 -- x"322D2C2F", x"2F2C2C30", x"2F2C2D30", x"312E2D2E", x"282B2E2E", x"2C2B2D30", x"2C2A2C2F", x"2D29282C",
									 -- x"2E2A292B", x"2C2A2A2C", x"2D2C2B2C", x"2F31302E", x"30303132", x"32323130", x"2D2E2E30", x"34323033",
									 -- x"33393937", x"3B3C3836", x"3737383A", x"3D3F3F3F", x"40414241", x"40424549", x"48494A4B", x"4C4B4A49",
									 -- x"4C4C4C4E", x"50515150", x"52525455", x"56585859", x"5858575A", x"5E5C5C61", x"60636565", x"66686765",
									 -- x"6567696A", x"6B6E7070", x"6F71716F", x"6E707273", x"7175746F", x"6E72726D", x"716F6E6E", x"6E6E6D6D",
									 -- x"6A686968", x"65686A67", x"65646362", x"61615F5E", x"5F5F5E5C", x"59585758", x"5D585A59", x"53545651",
									 -- x"4041403D", x"3B3B3C3C", x"3C3C3C3F", x"403E3A36", x"33312D2B", x"2B2D2A26", x"2D2B2928", x"28282828",
									 -- x"28262424", x"25242526", x"29262628", x"2B2B2B2A", x"2E303232", x"34373938", x"37393A39", x"393A3B3C",
									 -- x"3C3E4141", x"40404042", x"3D404243", x"4446494D", x"4F4F4F51", x"53555656", x"5D5C6061", x"5F666C69",
									 -- x"6E727376", x"79797A80", x"82888B8E", x"9496999F", x"A1A3A9B0", x"B4B6B9BA", x"C0C5C9CB", x"CACBCFD4",
									 -- x"D3D6DADB", x"DBDAD9D9", x"DBDDDEDD", x"DEE0E1E1", x"E0E2E3E3", x"E3E3E4E6", x"E5E4E6EA", x"EFF1F4F7",
									 -- x"F3F3F2F1", x"F0EDEAE7", x"E2E3E1E2", x"E7E9E9EC", x"EDEFF1F3", x"F4F5F8F9", x"F7F8FAFB", x"FDFDFDFD",
									 -- x"FEFEFFFF", x"FFFEFDFB", x"F8F7F7F7", x"F9F9F7F6", x"F5F6F6F4", x"F2F1F4F6", x"F5F3F0EF", x"EEEDEBE8",
									 -- x"E2DFDDDC", x"DBDADADB", x"DFE0E2E4", x"E6E8EBEC", x"EAEBEBEB", x"EBECECEC", x"EAEAE9E9", x"E9E8E6E3",
									 -- x"E1E3E4E6", x"E6E5E4E3", x"E6E5E3E0", x"E0E1E0DE", x"E0E0DDD9", x"D6D5D4D1", x"D0D1D2D1", x"D0D1D1CF",
									 -- x"CECECDCC", x"CCCCCBC9", x"C7C5C5C8", x"C8C6C5C7", x"C6C4C1BF", x"BFBFBEBD", x"BEBDBBBA", x"B8B7B5B3",
									 -- x"AFADAAA9", x"A9A8A6A4", x"A1A2A2A1", x"9F9E9D9E", x"9E9F9C9C", x"9F9E9B9C", x"9C9C9C9C", x"9B9A9999",
									 -- x"93929191", x"908E8B88", x"86858382", x"7F7B7979", x"79777777", x"76737273", x"7475777A", x"7B7B7B7B",
									 -- x"79797877", x"76757473", x"7271706D", x"6B696765", x"6262605E", x"5B595756", x"57555353", x"52514D4A",
									 -- x"4C4B4948", x"47474747", x"3E3F3F3E", x"3E3F3D3B", x"3B393737", x"38383430", x"32333434", x"32303031",
									 -- x"2F2B2C32", x"332F2D30", x"2E2B2C2F", x"2F2B2A2B", x"282B2E2E", x"2C2B2C2D", x"312E2D2C", x"29252629",
									 -- x"2E29272B", x"2F2D2B2B", x"29292B2C", x"2C2D2F31", x"30303132", x"32333334", x"30302E30", x"33323034",
									 -- x"363B3936", x"39393634", x"37383939", x"393B3E3F", x"3D3E3F3F", x"3E404347", x"47484949", x"48474849",
									 -- x"4B4A4A4B", x"4E4F4E4D", x"4F505153", x"54555656", x"5657575A", x"5E5B5A5F", x"61636566", x"66676665",
									 -- x"66686969", x"696B6C6C", x"6D6D6B6B", x"6D717372", x"6D6D6D6D", x"6C6B6A69", x"6D6C6C6A", x"6B6C6E6E",
									 -- x"67666766", x"63656763", x"62616060", x"605E5D5C", x"5A5C5E5C", x"58555759", x"5A555656", x"52535753",
									 -- x"3D3F3F3C", x"3B3B3C3C", x"3E3B3A3B", x"3C3B3938", x"32322F2B", x"292A2926", x"28272729", x"29272525",
									 -- x"26232223", x"24242425", x"24232427", x"2A2B2B2C", x"2E303131", x"32343534", x"37383939", x"3A3C3C3B",
									 -- x"3F404141", x"41414142", x"41434545", x"4546494C", x"504F4F51", x"54565656", x"5C5E6261", x"5F646968",
									 -- x"6C707174", x"7878797E", x"8086898C", x"9194989E", x"A3A3AAB1", x"B1B4B7B7", x"BEC2C6C8", x"C7C9CCD0",
									 -- x"D3D7DCDF", x"DEDDDCDC", x"DBDEDFDE", x"DEE0E1E1", x"E0E1E2E2", x"E1E1E2E3", x"E2E1E2E6", x"EAEDF0F4",
									 -- x"F4F4F4F4", x"F4F1EDEA", x"E7E7E2E1", x"E6E7E6E7", x"E6E9ECEE", x"EFF0F3F5", x"F3F5F7FA", x"FBFCFCFB",
									 -- x"FDFDFEFF", x"FFFFFEFD", x"FCFBFBFA", x"F9F7F5F4", x"F2F1F0EF", x"EEEFF2F5", x"F8F7F4F0", x"EEEEEDEB",
									 -- x"E3E2E0DF", x"DEDCDAD9", x"DFE0E0E1", x"E2E4E7E8", x"E8EAECEB", x"EAEBEBEB", x"E9EAEBEC", x"EDEDEAE6",
									 -- x"E4E4E3E3", x"E3E3E4E4", x"E2E1E0DF", x"E0E2E1DE", x"DEDFDEDA", x"D8D6D4D1", x"D1D3D3D2", x"D1D2D1CF",
									 -- x"CCCBCAC8", x"C8C8C8C6", x"C5C4C4C4", x"C4C3C3C3", x"C1C0BDBB", x"BBBCBBB9", x"B8B7B6B4", x"B3B2B0AF",
									 -- x"AAA9A7A6", x"A5A4A3A2", x"9D9D9E9E", x"9D9C9B9B", x"9A9A9798", x"9D9C999A", x"99999897", x"96959494",
									 -- x"918F8E8D", x"8C8A8684", x"84838280", x"7C777575", x"77757475", x"73707174", x"73747677", x"78787877",
									 -- x"75767573", x"71706E6C", x"6B6B6966", x"65656462", x"5D5C5B59", x"58565453", x"56524E4D", x"4E4E4B48",
									 -- x"48474543", x"41403F3F", x"3B3C3C3B", x"3B3B3A37", x"37363434", x"3536322E", x"30303132", x"312F2E2F",
									 -- x"2E2C2E32", x"33302D2D", x"2E2D2D2E", x"2D2B292A", x"282A2C2C", x"2C2B2B2B", x"302F2D2A", x"29282A2B",
									 -- x"2B28272A", x"2F302E2C", x"292B2E2E", x"2C2B3035", x"2F303032", x"33353636", x"32333130", x"33343335",
									 -- x"36393634", x"36363434", x"37393A38", x"383A3C3E", x"393B3F41", x"41424344", x"44454747", x"46464749",
									 -- x"4949494A", x"4C4D4C4B", x"4E4F5051", x"52535354", x"54575759", x"5C5A595D", x"62636465", x"66666665",
									 -- x"66686867", x"66676766", x"6A696767", x"6B6F706E", x"6866666A", x"6A666567", x"67686866", x"66686A6A",
									 -- x"66656664", x"6162635E", x"5D5C5C5D", x"5D5B5959", x"565B5E5D", x"59555556", x"55535455", x"53535350",
									 -- x"3D3F3F3D", x"3B3B3B3B", x"3C393839", x"39383738", x"3233312C", x"2A2C2B29", x"2928282A", x"2A272525",
									 -- x"27242224", x"26262524", x"23222326", x"27282A2D", x"2C2D2E2D", x"2E303130", x"35363637", x"3A3D3D3A",
									 -- x"403F3F40", x"42444444", x"47484848", x"494A4D4F", x"51525355", x"585A5B5B", x"59606260", x"62656667",
									 -- x"6A6D6D71", x"7676777D", x"7D84878B", x"9194979D", x"A2A1A8AF", x"ADAFB5B4", x"BABEC2C4", x"C5C7CACD",
									 -- x"D0D5DADD", x"DEDFE1E2", x"E1E2E3E2", x"E2E3E3E1", x"E1E2E2E2", x"E1E1E1E1", x"E0DFE1E3", x"E6E7EAED",
									 -- x"F1F1F1F3", x"F4F4F1EE", x"EDEBE4E1", x"E4E4E2E3", x"E2E4E7E9", x"EBECEDEE", x"EFF0F2F5", x"F6F7F8F8",
									 -- x"FAFAFAFC", x"FDFDFDFD", x"FDFDFBFA", x"F9F7F5F3", x"F0EEECEC", x"ECEBECEF", x"F4F5F3EF", x"EBEBEBEA",
									 -- x"E5E4E2E0", x"DFDEDCD9", x"DCDDDEDF", x"E0E1E3E5", x"E7E9EAE9", x"E9EBEAE8", x"E9EAEBEC", x"EDEFEDE9",
									 -- x"E7E6E4E3", x"E2E2E3E3", x"E0E1E1DF", x"DFE0DFDE", x"DEDFDEDC", x"D9D8D6D3", x"D3D4D4D3", x"D2D1D0CE",
									 -- x"CACBC9C6", x"C6C7C6C4", x"C5C7C6C2", x"C1C2C2C0", x"BDBDBAB7", x"B7B8B7B4", x"B3B1B0AE", x"ADACABAA",
									 -- x"A7A7A6A3", x"A09E9E9E", x"99999A9A", x"99989796", x"96959394", x"97969396", x"93939190", x"8F8E8D8D",
									 -- x"8C8B8988", x"88868380", x"817E7C7B", x"79757373", x"73707072", x"716D6E72", x"71717374", x"74747473",
									 -- x"6F71706D", x"6B6A6866", x"6665625F", x"5E5F5E5C", x"59575555", x"5553514E", x"504D4A49", x"4A4A4948",
									 -- x"4443413F", x"3C3B3B3B", x"3B3B3A37", x"37373633", x"32333230", x"3031312F", x"302E2D2F", x"2F2D2C2C",
									 -- x"2D2D2E2F", x"2F2E2D2C", x"2D2E2F2D", x"2C2C2A29", x"2A292929", x"2A2A2B2B", x"2C2D2C2A", x"2B2E2F2C",
									 -- x"28292829", x"2B2E2E2C", x"2D2F3130", x"2D2C3138", x"33333335", x"37383838", x"35383632", x"35363535",
									 -- x"36363333", x"35333133", x"35373837", x"37393A39", x"37393C3E", x"40404040", x"3F404243", x"44444444",
									 -- x"4747484A", x"4B4C4C4B", x"4C4D4D4E", x"4F505051", x"51565654", x"5758595B", x"5F606264", x"65666565",
									 -- x"63656665", x"65656564", x"66666565", x"676A6A69", x"67646367", x"66636265", x"62636362", x"63656360",
									 -- x"6161625F", x"5C5E5F5A", x"5958595B", x"5A585758", x"56585B5B", x"59565454", x"51525151", x"53514E4E",
									 -- x"3F41413E", x"3B3A3A39", x"3B393A3C", x"3D3A3839", x"3334322D", x"2C2F2F2C", x"302C2A2A", x"29272728",
									 -- x"2A272527", x"28272524", x"25242424", x"2525282B", x"292A2A29", x"2A2E3030", x"32323334", x"393D3C38",
									 -- x"3F3E3D40", x"44474847", x"49494949", x"4A4D5053", x"5355585B", x"5C5D6062", x"5760615F", x"64666465",
									 -- x"6B6D6C6F", x"7577797E", x"7C83878C", x"9295989D", x"9F9DA5AC", x"A9ACB3B3", x"B6B9BDC1", x"C4C7CACC",
									 -- x"CCD1D6DA", x"DCDFE4E8", x"E9E9E8E7", x"E9EAE7E3", x"E2E2E1E1", x"E1E1E0E0", x"E0DFE0E2", x"E3E4E6E8",
									 -- x"EAEAEAED", x"F0F2F1EF", x"EEEBE2DE", x"E1E0DDDD", x"DFDFE0E3", x"E6E8E7E6", x"EBECEEEF", x"F1F3F4F5",
									 -- x"F6F6F7F8", x"FAFBFBFB", x"FAF9F7F6", x"F6F5F3F1", x"F2EFEEEE", x"EDEBE9EA", x"EEF0F0EB", x"E8E7E8E7",
									 -- x"E6E5E3E1", x"E0DFDDDB", x"D8DADCDE", x"DEDFE1E2", x"E5E7E7E7", x"E9EAE8E5", x"E8E9E7E6", x"E8EBECEA",
									 -- x"E8E8E7E5", x"E4E3E2E1", x"E0E3E4E1", x"DEDDDDDC", x"DFE0DFDD", x"DBDAD8D6", x"D2D3D3D1", x"CFCECCCA",
									 -- x"CCCDCCC9", x"C9CAC8C5", x"C4C7C6C0", x"BEC1C0BC", x"BCBCB9B5", x"B4B4B2AF", x"AFAEACAA", x"A9A8A7A6",
									 -- x"A4A4A3A0", x"9B989798", x"96959494", x"9492908E", x"92929090", x"918E8D91", x"8E8D8C8A", x"89898888",
									 -- x"87858484", x"8483807E", x"7E7A7777", x"77757271", x"6E6C6D70", x"6E6A6B6F", x"6D6D6E6F", x"6F6F6F6E",
									 -- x"6B6D6C69", x"66666563", x"64635F5B", x"595A5956", x"55524F4E", x"4F4E4A47", x"4A494847", x"46444342",
									 -- x"4241403D", x"3B3A3B3B", x"38383633", x"3232312E", x"2E30302D", x"2A2B2E2F", x"312D2B2C", x"2C2A292A",
									 -- x"2C2C2C2A", x"2B2D2D2B", x"2A2D2E2B", x"292A2926", x"2B292727", x"282A2B2B", x"2A2E2E2A", x"2B302E28",
									 -- x"282B2B28", x"272B2D2C", x"2F2F302F", x"2C2B3037", x"39383839", x"3A3B3938", x"393E3A34", x"36383532",
									 -- x"36343132", x"34302D31", x"33343434", x"36383734", x"36353637", x"393A3A3A", x"3C3C3D3F", x"4243403E",
									 -- x"4546484A", x"4B4B4C4C", x"4949494A", x"4A4B4C4C", x"4E54534F", x"5256575A", x"5D5E6063", x"65656565",
									 -- x"63656766", x"65656462", x"64656564", x"64656665", x"68656464", x"62616162", x"62626161", x"6464605A",
									 -- x"5C5C5D5A", x"575B5D58", x"5757585A", x"59575658", x"58575656", x"57575655", x"4F524E4C", x"514F4B4E",
									 -- x"4242413F", x"3B373635", x"36373A3A", x"393C3B34", x"3434322F", x"2E2F2D2B", x"322D2A2B", x"2A272628",
									 -- x"25262728", x"28272422", x"21232527", x"27272627", x"29272628", x"2C2E2E2D", x"31303133", x"3637393B",
									 -- x"3B3D3F41", x"4244474A", x"464C4C4B", x"50505158", x"56585A5D", x"60616161", x"63626263", x"65656563",
									 -- x"656D7372", x"71757C7F", x"82838689", x"8E93989A", x"9BA0A4A5", x"A6AAAFB1", x"B3B5BBC1", x"C3C4C6C9",
									 -- x"CBCED2D8", x"DCDEE1E4", x"E8E9E6E7", x"EBECECEE", x"EBEAE9E8", x"E6E5E2E1", x"E2E2E2E2", x"E2E3E4E6",
									 -- x"E7E6E5E6", x"E8EAEBEA", x"E8E4E0DF", x"DEDCDBDC", x"DBDDDFE0", x"E1E1E3E4", x"EAECEDEE", x"EEEFF1F2",
									 -- x"F3F3F4F7", x"F7F5F6F8", x"F7F7F5F4", x"F2F1F0F0", x"F0EFEFEE", x"EDECEAEA", x"EBEDEDE9", x"E7E8E6E2",
									 -- x"E6E7E3DB", x"D8DADAD6", x"D5D7D9DA", x"DADADDDF", x"DFE1E2E4", x"E6E6E5E4", x"E3E3E3E4", x"E6E7E7E7",
									 -- x"E7E5E4E5", x"E5E3E2E3", x"E2E4E4E3", x"E1DFDEDD", x"DDDDDCDC", x"DBD9D7D5", x"D5D4D2D0", x"CECDCCCB",
									 -- x"CBCBCAC8", x"C5C5C6C8", x"C6C4C2C2", x"C3C2BFBB", x"BAB8B7B6", x"B2AFAFB2", x"ABA9A7A6", x"A7A7A5A3",
									 -- x"9F9C9A9A", x"98959495", x"97959290", x"90908F8E", x"8C8D8E8D", x"8C8C8A88", x"86898986", x"85868480",
									 -- x"80807F7F", x"7F7D7B79", x"7B767374", x"74716D6C", x"6B6C6A65", x"64686967", x"6968686A", x"6C6C6966",
									 -- x"68676562", x"6262605D", x"5D5B5856", x"55555555", x"4F4E4C4B", x"4B4B4A49", x"46444241", x"41413F3E",
									 -- x"3A3E3E3A", x"38393835", x"37333133", x"33312D2C", x"2F2F2E2D", x"2C2C2E2F", x"2B2D2E2B", x"28282928",
									 -- x"2B2C2D2D", x"2C2C2C2C", x"2D2C2B2A", x"2A2B2A2A", x"28282829", x"2A2B2928", x"282A2B2B", x"2A292A2C",
									 -- x"2E2A282A", x"2A292A2E", x"2E2C2E33", x"3230333A", x"3A39393A", x"3938393B", x"3E3E3D3B", x"3A3B3A38",
									 -- x"37373533", x"3233322F", x"34333232", x"33343332", x"3536343C", x"383D3C40", x"3B3D3E3D", x"3F414240",
									 -- x"40434546", x"47494846", x"4748494B", x"4D4D4D4C", x"4B4E5050", x"4E50555A", x"545C6160", x"60636462",
									 -- x"64605F61", x"63616062", x"60606264", x"63606061", x"6261605D", x"5B5B5C5C", x"5F605F5C", x"5A595857",
									 -- x"5B5C5A57", x"585B5B57", x"58565554", x"54555555", x"53525356", x"5754504D", x"4F4F4E4F", x"53504C4D",
									 -- x"42413E3B", x"3837383A", x"35363837", x"35383730", x"30302F2D", x"2D2D2C2A", x"2F2B2A2C", x"2C292729",
									 -- x"27272727", x"27272726", x"26252423", x"24262829", x"2A282627", x"2A2D2E2F", x"2F2E2F32", x"3435383B",
									 -- x"3B3B3B3C", x"3F424546", x"4B4D4E4F", x"5355575A", x"58595B5E", x"60626262", x"64636262", x"63646667",
									 -- x"686C6E6E", x"6D71787C", x"7F7F8184", x"8A909698", x"9A9B9B9D", x"A3AAADAC", x"B3B3B6BB", x"BEC0C1C3",
									 -- x"C8CACED3", x"D6D9DDE1", x"E4E6E5E6", x"ECEEEEF1", x"F1F0EFEE", x"EEEDECEB", x"E9EAEAE9", x"E8E6E6E5",
									 -- x"E9E8E7E7", x"E7E8E7E6", x"E3E1E0E0", x"DFDCDAD9", x"DADCDDDE", x"DFDFE1E2", x"E7E8EAEC", x"ECEDEFF0",
									 -- x"F1EFEEEF", x"F0F0F3F7", x"F5F4F3F2", x"F0EEEDEC", x"EBECEDED", x"EDEBEAE9", x"EAECECE8", x"E6E7E6E2",
									 -- x"E3E4E1DB", x"D9D9D8D5", x"D3D4D5D6", x"D7D8D9D9", x"DBDEE0E1", x"E1E1E1E2", x"E2E1E1E2", x"E3E3E3E2",
									 -- x"E4E2E2E4", x"E4E2E2E2", x"DFE0E0DF", x"DDDBDBDC", x"DDDDDCDB", x"DAD8D5D3", x"D3D3D2D0", x"CECCCAC9",
									 -- x"C8C8C8C7", x"C7C6C4C3", x"C3C2C2C2", x"C2C0BBB7", x"BAB6B4B4", x"B3B0AEAD", x"A8A6A5A4", x"A4A4A3A2",
									 -- x"9D9A9898", x"97949292", x"9392908F", x"8F8F8F8E", x"898A8988", x"88898785", x"82838381", x"807F7E7C",
									 -- x"7A7A7A78", x"76757575", x"75727071", x"716D6866", x"66686763", x"63666764", x"63656767", x"64626263",
									 -- x"6162615E", x"5D5C5B59", x"58565452", x"5150504F", x"4A4A4A48", x"47464646", x"4342403F", x"3E3D3C3B",
									 -- x"3A3C3C38", x"36373532", x"32303031", x"312E2D2E", x"2E2D2C2B", x"2A292A2B", x"292A2A2B", x"2A292929",
									 -- x"28292A2B", x"2A2A2A2A", x"2C2B2A29", x"2A2B2B2B", x"28272627", x"27272725", x"2426292A", x"29282829",
									 -- x"2C28282C", x"2F2D2C2D", x"2A2A2C31", x"35363A3E", x"3A38383A", x"3B3A3A3B", x"42424240", x"3F3E3C3A",
									 -- x"38353334", x"34302F30", x"31303031", x"33343333", x"33333338", x"383B3A3D", x"3B3D3D3D", x"3E414241",
									 -- x"40414140", x"41444646", x"46464648", x"494A4A49", x"46494B4C", x"4B4D5256", x"5156595A", x"5B5D5E5E",
									 -- x"5E5E5F5F", x"5D5B5C5E", x"5D5D5F62", x"62605E5E", x"5E5E5C5A", x"595A5B5C", x"58585858", x"57565657",
									 -- x"55575755", x"56595956", x"58565453", x"53535354", x"52504F51", x"52504D4C", x"52514E4F", x"514F4C4E",
									 -- x"403F3C3A", x"38393B3D", x"3B3A3B3A", x"373A3A35", x"30312F2D", x"2D2E2D2A", x"2E2B2A2B", x"2B29282A",
									 -- x"2A2A2928", x"2829292A", x"2A272423", x"2527292A", x"28272625", x"27292C2E", x"2D2D2F31", x"3233363A",
									 -- x"3C3B3A3B", x"3F424546", x"4C4B4E52", x"55595C5B", x"5B5C5E61", x"63646464", x"65656564", x"6566686A",
									 -- x"69686A6D", x"7073787C", x"7D7C7D80", x"868D9296", x"9C9B999A", x"9FA5A7A6", x"B1B0B2B7", x"BCBFC1C3",
									 -- x"C6C7CACE", x"D1D4D8DD", x"DFE2E2E5", x"EBEEEEF0", x"F4F3F2F2", x"F2F2F2F1", x"F0F1F2F2", x"EFECE9E8",
									 -- x"E8E7E6E6", x"E7E7E6E5", x"E0DFDFE0", x"DEDAD9D9", x"DADBDCDD", x"DDDDDFE0", x"E3E5E7E9", x"EAEBECEC",
									 -- x"EFEDECEC", x"ECEDF1F4", x"F4F4F4F4", x"F2EFEDEB", x"EAEBEBEB", x"EBEAEBEB", x"EBECEBE8", x"E6E7E6E4",
									 -- x"E0DFDEDC", x"D9D7D5D3", x"D1D0D0D1", x"D2D4D3D3", x"D6D9DCDC", x"DBDADCDE", x"DFDFE0E1", x"E2E2E1E0",
									 -- x"E0DFDEE0", x"E0DFDEDE", x"DEDEDDDC", x"DADADBDC", x"DCDBD9D8", x"D6D4D2D1", x"D0D0D0CF", x"CDCBC9C7",
									 -- x"C5C4C3C3", x"C5C4C2C0", x"C1C1C0C0", x"BFBDB9B7", x"B8B4B1B2", x"B3B1ACA8", x"A9A7A5A2", x"9F9D9B9B",
									 -- x"9B989595", x"9593908F", x"8D8D8D8D", x"8C8C8C8C", x"89888685", x"86878683", x"817F7F7F", x"7E7B797A",
									 -- x"76777674", x"706F7173", x"716F6F70", x"706C6764", x"63666664", x"64656461", x"61636462", x"5F5D5D5E",
									 -- x"5D5E5E5B", x"59595856", x"5352504E", x"4D4C4A4A", x"46474745", x"42404142", x"3E3E3E3C", x"3B393838",
									 -- x"37383734", x"3334322F", x"2D2E2E2F", x"2D2C2C2D", x"2C2C2B2A", x"29282929", x"2927272A", x"2B292829",
									 -- x"28292A2B", x"2B2A2A2A", x"29282726", x"27282828", x"28272525", x"24242423", x"24252626", x"25252728",
									 -- x"2A26262B", x"2F2F2E2E", x"2D2C2D31", x"363A3B3C", x"3D3B3B3E", x"403F3E3E", x"41424241", x"41403E3B",
									 -- x"39343336", x"352F2D30", x"2F2F3031", x"32333232", x"34323334", x"39373938", x"393A3A3A", x"3B3D3E3E",
									 -- x"40403F3E", x"3E414343", x"42424243", x"45474747", x"47484949", x"48494A4C", x"50505256", x"5757595B",
									 -- x"5A5B5B5A", x"5A5B5B5A", x"5C5B5B5E", x"5F5D5B5A", x"5C5B5A59", x"57565758", x"54535355", x"55535356",
									 -- x"54565653", x"52545452", x"56545250", x"4F4F5050", x"514E4C4D", x"4D4C4C4C", x"504F4B4B", x"4D4B494C",
									 -- x"3D3D3E3E", x"3D3D3D3D", x"3A393A38", x"36393A36", x"35353432", x"31312F2C", x"312D2B2A", x"2928292B",
									 -- x"2D2D2D2C", x"2C2C2C2C", x"2B292728", x"292A2928", x"27272726", x"26282B2E", x"2D2D3032", x"32323438",
									 -- x"3A3A3B3D", x"3F434648", x"4A484E54", x"555A605D", x"60616466", x"6768696A", x"696A6A6C", x"6D6D6D6C",
									 -- x"6D6B6C73", x"7778797B", x"7C7D7F81", x"84898F93", x"9B9C9E9E", x"9EA0A5A8", x"AEAEB0B5", x"B8BBBDC0",
									 -- x"C5C5C8CB", x"CED1D6DB", x"DBDFE0E2", x"E8E9E9EB", x"F1EFEEED", x"EDECECEC", x"EEEFF2F2", x"F1EEECEB",
									 -- x"E7E6E6E6", x"E6E5E5E4", x"E2E1E0DF", x"DCD9D9DB", x"DCDBDBDB", x"DBDCDDDD", x"E0E2E4E6", x"E7E8E8E8",
									 -- x"EAEBECEC", x"ECECEDEE", x"F2F3F4F4", x"F3F0EDEB", x"EBEAE9E7", x"E6E7E9EC", x"EAEBEAE7", x"E5E5E4E2",
									 -- x"DDDBDBDA", x"D8D5D3D3", x"CFCFCFCF", x"CFCFCFCF", x"D2D4D5D5", x"D5D5D7D8", x"DADADCDE", x"DFE0DFDE",
									 -- x"DDDCDBDB", x"DBDAD9D8", x"DBDADAD9", x"D9D9DADA", x"DAD8D7D5", x"D4D2D0CF", x"CDCDCDCC", x"CBC9C8C7",
									 -- x"C4C2C0BF", x"BFC0C0C0", x"C0BFBDBC", x"BABABABA", x"B7B3B0B0", x"B1AFAAA6", x"A9A7A5A2", x"9E999696",
									 -- x"98969393", x"93928F8D", x"88898B8A", x"88878788", x"87868483", x"8485837F", x"817D7C7F", x"7D787679",
									 -- x"75757472", x"6F6E6F71", x"6D6D6D6E", x"6F6C6865", x"62646462", x"61615F5D", x"615E5C5C", x"5D5D5B58",
									 -- x"5A5A5957", x"57575552", x"4E4D4B4A", x"49474544", x"45454442", x"403E3D3C", x"393A3B3A", x"38363637",
									 -- x"33343331", x"3133322F", x"2C2C2C2C", x"2B2A2A2A", x"2A2A2A2A", x"29292A2B", x"2925252A", x"2C282628",
									 -- x"292A2B2B", x"2A2A2A2B", x"27272626", x"26252524", x"28262523", x"22222323", x"27262523", x"22232527",
									 -- x"29252427", x"2A2C2D2F", x"302F2E30", x"353A3A37", x"3E3D3E40", x"41403F40", x"3C3D3E3E", x"3E3F3E3B",
									 -- x"3A373638", x"36322F2F", x"31313232", x"32323131", x"37333531", x"38343734", x"39393838", x"393A3B3C",
									 -- x"3E3F4040", x"40403F3E", x"403F3F40", x"43454647", x"47474848", x"48484848", x"4D4C4E52", x"52505359",
									 -- x"57565453", x"575C5B55", x"5B58585A", x"5B595756", x"57575757", x"56545455", x"57545456", x"54505053",
									 -- x"54565552", x"50505151", x"51504F4D", x"4C4C4D4E", x"504D4B4B", x"4C4B4C4D", x"4B4A4849", x"4C4A4749",
									 -- x"3E3F4042", x"42413F3E", x"3B3A3A3A", x"37393B39", x"38383735", x"34343230", x"312F2E2D", x"2C2B2B2C",
									 -- x"2F313233", x"32302F2E", x"2C2B2A2B", x"2D2D2A28", x"28292A2A", x"29292B2D", x"2C2D3034", x"34343537",
									 -- x"35383C3E", x"40424649", x"4A495156", x"555B6261", x"6466696B", x"6C6D6F70", x"72717173", x"76767472",
									 -- x"78747478", x"7B797879", x"7D818586", x"86878C91", x"97999C9F", x"A0A3A6A9", x"A9ABAFB2", x"B2B2B5B9",
									 -- x"C4C4C6CA", x"CCCFD4D8", x"D8DCDDDF", x"E4E4E3E6", x"EAE9E7E5", x"E4E3E2E1", x"E5E7E9EA", x"EAE9E9E8",
									 -- x"E6E6E5E4", x"E3E3E3E3", x"E4E3E3E3", x"DFDCDBDC", x"DCDCDBDA", x"DADADADB", x"DBDDDFE1", x"E3E4E4E4",
									 -- x"E4E6E8E9", x"E9E9E9E9", x"ECEDEFF0", x"EFEDEBE9", x"E9E9E8E5", x"E3E3E4E6", x"E8E8E7E4", x"E3E2E0DE",
									 -- x"DCDAD9D8", x"D6D3D2D3", x"CFD0D1CF", x"CDCCCDCE", x"D0CFCECF", x"D1D3D3D2", x"D3D4D5D8", x"DADADAD9",
									 -- x"D9D9D8D7", x"D7D7D6D4", x"D5D5D5D5", x"D6D6D6D6", x"D7D6D5D4", x"D3D2D0CF", x"CCCCCBC9", x"C8C7C6C6",
									 -- x"C3C3C1BE", x"BCBBBBBC", x"BCBBBAB8", x"B8B8B9B9", x"B5B3B0AE", x"ADACA9A6", x"A4A3A2A2", x"9E999798",
									 -- x"96949290", x"91918F8C", x"87898989", x"86848484", x"83838280", x"81807D79", x"7D78777A", x"79737276",
									 -- x"7271706E", x"6D6C6B6B", x"6A6A6969", x"68676462", x"5F605F5E", x"5C5B5A58", x"5A585656", x"58595755",
									 -- x"56555452", x"5354514D", x"49484746", x"45434140", x"42403E3E", x"3E3D3A38", x"36383938", x"36353536",
									 -- x"32323130", x"3030302E", x"2C2B2929", x"2A2B2A28", x"29292A2A", x"2A29292A", x"2824242A", x"2C282628",
									 -- x"2A2A2928", x"27272829", x"29282828", x"28262422", x"25242321", x"20202122", x"24242322", x"21222324",
									 -- x"25252526", x"27282B2E", x"2D2C2B2E", x"34393A37", x"393A3C3E", x"3C3A3B3D", x"3B3C3C3C", x"3D3F3F3D",
									 -- x"3B3D3C38", x"3636332F", x"33333333", x"32323231", x"3733352F", x"35313533", x"3B3A3939", x"39393A3B",
									 -- x"3B3C3D3F", x"403E3D3D", x"403F3E3F", x"41434445", x"42424445", x"47494949", x"49484A4E", x"4C494D55",
									 -- x"51514F4D", x"50555552", x"58555355", x"56565454", x"50505255", x"55535254", x"55535253", x"524E4E51",
									 -- x"4F51504E", x"4D4E5152", x"4E4D4D4B", x"4A4A4C4E", x"4C4A4A4B", x"4B4B4B4C", x"4749494B", x"4F4D494A",
									 -- x"43434243", x"43434241", x"403E3E3E", x"3A3B3D3C", x"393A3938", x"37373633", x"2F313333", x"32302F2E",
									 -- x"32343738", x"37353333", x"302F2E2E", x"2E2F2E2D", x"2A2B2D2D", x"2C2B2B2C", x"2C2D3034", x"36363637",
									 -- x"34393F42", x"4244484D", x"494B5155", x"55595F61", x"65686B6D", x"6E707375", x"7B7A7879", x"7B7D7D7C",
									 -- x"7F7D7B7C", x"7C7C7D7F", x"82878C8D", x"8B8B8E92", x"9B98989D", x"A3A5A3A1", x"A3A6ABAE", x"AFAFB4BA",
									 -- x"C1C1C4C7", x"CACBCFD4", x"D3D8D9DB", x"DFE0E0E3", x"E5E4E2E0", x"DFDEDCDB", x"DEDFE0E1", x"E1E1E1E2",
									 -- x"DFE0E0E0", x"E1E2E4E5", x"E4E4E7E8", x"E6E1DEDD", x"DEDDDCDB", x"DBDADAD9", x"D8D9DADD", x"DFE1E1E0",
									 -- x"E0E2E3E4", x"E5E7E9E9", x"E7E8EAEB", x"EBEAE9E8", x"E7E9EAE9", x"E5E3E2E2", x"E7E7E7E5", x"E3E1E0DE",
									 -- x"DBDBD9D7", x"D5D4D3D3", x"D0D1D2D0", x"CCCACBCD", x"CDCBCACB", x"CED0CFCD", x"D0D0D1D3", x"D4D5D4D3",
									 -- x"D4D5D4D4", x"D4D5D4D3", x"D2D1D1D2", x"D3D3D3D2", x"D4D3D2D2", x"D2D1D0CF", x"CDCCCAC8", x"C6C4C4C3",
									 -- x"C2C3C3C1", x"BCB9B8B8", x"B8B8B8B8", x"B8B7B5B4", x"B4B3B0AC", x"A9A8A7A6", x"A3A1A0A0", x"9D989595",
									 -- x"9392908E", x"8D8D8C8B", x"87888887", x"85848382", x"8182817F", x"7D7C7976", x"78747375", x"74706F72",
									 -- x"6F6E6C6C", x"6B6A6866", x"67676663", x"6262605E", x"5C5C5C5B", x"5A595857", x"53555655", x"53535557",
									 -- x"52525150", x"50504D49", x"48474544", x"4442403F", x"3C3A3839", x"3B3B3835", x"35353635", x"34333333",
									 -- x"3131312F", x"2D2C2C2C", x"2A292727", x"2A2C2B28", x"28292A29", x"28272727", x"26242529", x"2B29292A",
									 -- x"2B2B2A29", x"27272828", x"27272728", x"27262321", x"2221201F", x"1E1E1F20", x"1D1E2022", x"23222121",
									 -- x"22252829", x"2928292B", x"2B2A2A2D", x"31343636", x"35373A3B", x"3836373B", x"3F403F3E", x"3E403F3E",
									 -- x"3B3E3D37", x"3538352F", x"33333333", x"32333334", x"3232322F", x"31313433", x"38373737", x"37373739",
									 -- x"38373739", x"3A3B3D3F", x"3F3E3D3D", x"3F404141", x"3F3F4142", x"43444546", x"4747494C", x"4A474A50",
									 -- x"4B4F504D", x"4A4B4F52", x"52504F50", x"52525152", x"504F5053", x"524E4D4F", x"4C4D4D4D", x"4D4D4D4E",
									 -- x"4D4D4C4A", x"494B4C4E", x"4B4C4C4B", x"4A4B4C4E", x"48474849", x"49484849", x"4647484B", x"4F4C4849",
									 -- x"46454444", x"45444342", x"3F3D3E3E", x"3A3A3D3C", x"3D3E3E3C", x"3C3C3A37", x"34363737", x"35343332",
									 -- x"35383A3A", x"3938393A", x"36353534", x"34343435", x"2F303131", x"302F2E2D", x"302F2F33", x"36363636",
									 -- x"383C4043", x"44474B4E", x"4C4F5152", x"56595B5F", x"6366696C", x"6E707476", x"7D7E8080", x"80818385",
									 -- x"83858584", x"83858889", x"8A8D9294", x"94949597", x"A19D9CA0", x"A4A3A09D", x"A2A4A9AD", x"AFB1B7BD",
									 -- x"BDBEC1C5", x"C7C8CBCF", x"CDD2D4D6", x"DADBDCDF", x"E1E0DFDF", x"DFDEDDDC", x"DBDCDDDD", x"DDDDDDDE",
									 -- x"DADBDCDC", x"DDDFE3E5", x"E4E4E7EB", x"EBE7E3E1", x"E2E1E0DF", x"DFDEDCDA", x"DBDADADB", x"DDDDDDDC",
									 -- x"DDDFE0DF", x"E0E3E5E5", x"E5E6E7E7", x"E8E8E8E8", x"E6E8E9E8", x"E4E2E2E3", x"E5E5E6E5", x"E4E2E0DF",
									 -- x"DADCDBD6", x"D5D5D4D1", x"D0D1D0CE", x"CBC9C9C9", x"C9C8C8C9", x"CBCCCCCB", x"CDCDCECE", x"CFD0CFCE",
									 -- x"CFD0D0CF", x"CFD1D0CE", x"D0CECDCD", x"CFD0D0CF", x"CFCFCECE", x"CECDCCCA", x"CACAC9C7", x"C6C4C3C2",
									 -- x"C1C1C1C0", x"BEBCBAB9", x"BAB9B8B8", x"B8B7B3B0", x"B2B1AEA9", x"A7A7A6A3", x"A49F9C9C", x"99949191",
									 -- x"90918F8A", x"88888988", x"84848383", x"83828180", x"7F80807C", x"79777573", x"73717070", x"6F6D6D6E",
									 -- x"6B6B6A69", x"67656464", x"62636260", x"5F5F5E5B", x"5B5A5A5A", x"59575555", x"51535453", x"51505254",
									 -- x"4D50504E", x"4B4A4847", x"45444342", x"41403F3E", x"39373637", x"39383633", x"34343232", x"3131302F",
									 -- x"2F2F302D", x"2A28292B", x"28292826", x"282A2A28", x"27282929", x"28272626", x"25262729", x"292A2A2B",
									 -- x"292A2A2A", x"29282828", x"24242425", x"25252423", x"2121201E", x"1D1C1D1E", x"1C1D1F21", x"22232221",
									 -- x"23252728", x"29292929", x"2B292A2D", x"2F2E3034", x"36363839", x"3836383B", x"3E3F3F3D", x"3D3E3C3A",
									 -- x"393A3936", x"35363431", x"31323231", x"31323436", x"2F323232", x"2F323233", x"33323234", x"34333435",
									 -- x"35333334", x"36373A3E", x"3B3A3A3A", x"3C3D3E3E", x"3E3E3F3F", x"3E3E3F40", x"4847474A", x"4A49484A",
									 -- x"4A4A4C4C", x"4A494A4E", x"4D4C4D4E", x"4E4D4C4D", x"514E4E4F", x"4D49484B", x"474A4B49", x"494C4C4B",
									 -- x"4B4A4948", x"48484848", x"494A4B4B", x"4A4A4B4D", x"46454647", x"46444445", x"46464446", x"4A484547",
									 -- x"45454546", x"47464341", x"42404243", x"40404444", x"43444341", x"40403D3B", x"3C3C3A37", x"35353637",
									 -- x"383A3B3A", x"393A3D3F", x"393A3C3C", x"3B3A3939", x"37373736", x"36353333", x"35312F31", x"34353434",
									 -- x"3A3B3E40", x"43474A4D", x"52555253", x"5A5B5A5F", x"6063676A", x"6C6F7376", x"7A7F8586", x"84838588",
									 -- x"888E918E", x"8C8D8E8D", x"91939598", x"9B9C9D9C", x"A1A0A2A4", x"A4A2A2A4", x"A8A7A8AB", x"ADB0B5B9",
									 -- x"BBBCC0C4", x"C6C7C9CC", x"C9CECFD1", x"D5D6D7DB", x"DDDDDDDE", x"DFE0DFDE", x"DCDCDDDE", x"DDDDDDDE",
									 -- x"DDDDDCDA", x"D9DADDDF", x"E5E4E6E9", x"EBEAE8E7", x"E6E5E4E3", x"E3E1DFDD", x"E0DFDDDC", x"DCDBDAD8",
									 -- x"D9DCDDDC", x"DCDEDEDD", x"E4E4E4E4", x"E5E6E7E7", x"E5E5E4E1", x"DEDDE0E3", x"E0E1E2E3", x"E2DFDDDC",
									 -- x"DADDDCD7", x"D5D7D5D0", x"D1CFCECC", x"CBC9C7C6", x"C6C7C8C8", x"C9C9C9CA", x"C9C9C8C9", x"CACBCBCA",
									 -- x"CDCECDCB", x"CBCCCBC8", x"CCCAC8C8", x"C9CBCCCC", x"CACACACB", x"CAC9C7C5", x"C6C7C7C7", x"C7C5C4C3",
									 -- x"C1BFBDBC", x"BEBFBFBF", x"C0BDB9B7", x"B7B6B3B1", x"B1B0ACA8", x"A6A6A4A1", x"A19A9697", x"96939192",
									 -- x"8F908E88", x"84848586", x"81807F7F", x"8081807F", x"7C7E7D78", x"73717070", x"6E6D6C6B", x"6B6A6A6A",
									 -- x"67686865", x"62606062", x"5B5D5E5C", x"5C5D5C5A", x"59595959", x"57545150", x"514F4E4E", x"50504E4C",
									 -- x"474B4E4A", x"45424343", x"403F3D3D", x"3C3B3B3A", x"39383838", x"37363432", x"3432302F", x"2F2F2D2C",
									 -- x"2B2D2E2C", x"2826282B", x"282A2927", x"26272827", x"26272929", x"29282827", x"26292A29", x"28292A2A",
									 -- x"25272829", x"28272525", x"24242324", x"25272828", x"2122211F", x"1D1D1D1E", x"21201F1F", x"20222324",
									 -- x"25252425", x"26292929", x"2826292E", x"2E2C3036", x"36353637", x"3838393B", x"393B3B3A", x"3A3A3835",
									 -- x"38363435", x"35333233", x"31313130", x"2F303335", x"2E353436", x"2F343133", x"31303133", x"34333335",
									 -- x"34323234", x"3535373A", x"36353637", x"3A3B3D3D", x"3A3C3D3D", x"3C3C3E40", x"46444346", x"48484643",
									 -- x"49434247", x"4C4B4746", x"4B4B4D4E", x"4C494748", x"4D49494B", x"4A484A4F", x"474C4D48", x"474B4B48",
									 -- x"47464648", x"4A4A4948", x"46484A4A", x"4848494A", x"46454546", x"45424243", x"49474343", x"46444346",
									 -- x"474A4B4A", x"494A4B4B", x"4B494644", x"44454849", x"4A484644", x"42414040", x"3E3F3E3B", x"3B3E3E3B",
									 -- x"3D3E3E3E", x"3F40403F", x"3D404240", x"3E3D3E3D", x"413F3D3C", x"3A38383B", x"35343436", x"36363739",
									 -- x"373C4244", x"45474C50", x"545B5B59", x"5B5F6163", x"6465686D", x"7277797A", x"7F82878A", x"88878A8E",
									 -- x"8E8F9193", x"95959594", x"9C9C9EA1", x"A4A5A4A3", x"A9AAAAAA", x"ABADADAB", x"AEAFB1B2", x"B4B8BCC0",
									 -- x"BFC0C4C8", x"C9C7C5C6", x"C8CBCECF", x"CED1D6DB", x"DDE0DFDC", x"DEDEDEE0", x"DEDDDDDE", x"DFE0DEDD",
									 -- x"DEDFDFDE", x"DDDCDCDC", x"E2E4E5E4", x"E5E7E7E6", x"E9E7E6E6", x"E5E3DFDD", x"E1DEDCDB", x"DBDAD8D6",
									 -- x"D7D7D8DB", x"DCDBDCDD", x"E0E1E0E0", x"E2E5E5E3", x"E2E2E2E0", x"DEDDDEE0", x"DDDEDEDE", x"DDDDDCDC",
									 -- x"DDD9D8DB", x"DBD6D3D2", x"CFCFCDCB", x"CACBC8C3", x"C5C7C5C3", x"C4C7C7C4", x"C6C5C4C3", x"C4C4C5C5",
									 -- x"C6C5C6C7", x"C7C4C4C6", x"C5C7C9C8", x"C5C5C7CA", x"C8C8C8C8", x"C7C6C5C4", x"C1C1C0BF", x"BDBCBBBB",
									 -- x"B8B6B6B8", x"BABBBDC1", x"C3BFBBB9", x"B9B8B6B3", x"AEADABA7", x"A5A3A09C", x"98989696", x"9493908F",
									 -- x"8E8C8986", x"83828180", x"7E7E7E7E", x"7E7C7B79", x"78777575", x"74736F6D", x"6C6B6A69", x"68666463",
									 -- x"6464625F", x"5E5F605F", x"5E5C5856", x"57595653", x"51535454", x"53515050", x"504F4C49", x"494A4845",
									 -- x"49484645", x"4342403F", x"3F3D3C3C", x"39363537", x"35343332", x"33333333", x"2D2E2F30", x"2F2D2A27",
									 -- x"26292A29", x"292A2825", x"28282929", x"28262525", x"29252325", x"28292828", x"29282829", x"2A2B2927",
									 -- x"21272724", x"24242426", x"25242221", x"20202123", x"2223221F", x"1D1E1F1E", x"201D1B1C", x"1F21201F",
									 -- x"21222223", x"24252727", x"272C2A2B", x"312F2B31", x"31313335", x"34343639", x"3B393633", x"32313132",
									 -- x"3734312F", x"2F2E2E2F", x"2F313130", x"3235332D", x"33333331", x"2F303336", x"302C2D32", x"332F3035",
									 -- x"34313032", x"32313133", x"30343737", x"37393A39", x"3B38393E", x"403E3D3E", x"3E3F4042", x"43444444",
									 -- x"42414041", x"43454645", x"43454747", x"46454445", x"4B494646", x"47494847", x"49494745", x"45474847",
									 -- x"43444443", x"44474948", x"45454543", x"42434547", x"46484948", x"46444343", x"43454544", x"44464644",
									 -- x"4A4D4F4F", x"4E4E4D4B", x"504E4B48", x"47474849", x"49494949", x"49484646", x"45474642", x"4142423F",
									 -- x"41434342", x"43434240", x"40414241", x"41424241", x"42414244", x"423F3D3E", x"403D3B3A", x"3A393B3D",
									 -- x"3C3F4345", x"46494E52", x"565A5B5C", x"61646567", x"67686B70", x"75797A7A", x"7F83898D", x"8C8A8B8D",
									 -- x"8E919699", x"9A9B9C9D", x"9D9EA1A4", x"A8A9AAA9", x"B0B1B1B2", x"B4B6B5B2", x"B2B4B5B6", x"B8BBBEC1",
									 -- x"C4C4C7CA", x"CAC9C8CA", x"CACCCED1", x"D3D7DBDE", x"DFE4E5E5", x"E8E8E7E9", x"E9E7E5E4", x"E4E3E2E0",
									 -- x"DEE0E2E2", x"E1E0E1E2", x"DFE0E1E0", x"E1E3E4E3", x"E1E1E1E3", x"E4E4E2E0", x"DBDBDCDC", x"DBDAD8D7",
									 -- x"D7D6D6D7", x"D8D7D8DA", x"D9DCDEDF", x"E0E1E1DF", x"E1E1E1E0", x"DFDFE0E1", x"DCDDDEDE", x"DDDCDBDB",
									 -- x"DCDCDCDC", x"DCDBD8D4", x"CFCECAC7", x"C6C6C4C0", x"C3C2C1BF", x"BFC1C0BE", x"C0BFBEBE", x"BFC0C0C0",
									 -- x"C2C1C2C3", x"C3C1C2C4", x"C0C2C4C4", x"C2C1C2C4", x"C2C2C2C2", x"C2C2C1C1", x"BCBCBBBA", x"B8B7B7B7",
									 -- x"B6B4B3B6", x"B9BABBBD", x"BEBBB8B6", x"B5B4B1AE", x"A9A8A5A1", x"9F9E9A97", x"97969593", x"92908E8C",
									 -- x"87868482", x"8180807F", x"7C7C7B7B", x"79777674", x"7573716F", x"6F6D6A67", x"67666463", x"6261605F",
									 -- x"5E5F5F5C", x"5B5B5957", x"59585553", x"52535250", x"4F505151", x"4F4E4E4E", x"494A4947", x"47494948",
									 -- x"46454443", x"42403E3C", x"3C3A3A3B", x"3A363332", x"32323233", x"3332302F", x"2F2E2D2C", x"2C2D2C2C",
									 -- x"292A2926", x"25272827", x"25242425", x"27262523", x"27262729", x"2A292828", x"272A2C2B", x"27252527",
									 -- x"21252421", x"23242223", x"24232322", x"21202121", x"23242421", x"1F20201F", x"1E1D1C1D", x"1F21201F",
									 -- x"20212223", x"24242526", x"282B292A", x"2F2C292E", x"2E2E2F31", x"32313133", x"39373431", x"30303131",
									 -- x"31303030", x"30303031", x"2D2F2F2D", x"2F32322E", x"2E2F302E", x"2C2C2E30", x"2F2B292B", x"2C2C2F33",
									 -- x"32302F30", x"30303133", x"31343535", x"35363837", x"35353639", x"3B3A3A3B", x"3B3D3E3E", x"3C3C3D3F",
									 -- x"3E3E3F40", x"40404141", x"3E404243", x"43434344", x"45444343", x"45464543", x"45444241", x"42454644",
									 -- x"42434341", x"42444645", x"44444442", x"41404142", x"42434545", x"45444444", x"42454644", x"43444544",
									 -- x"4C4E4F4F", x"50504F4C", x"4E4D4C4C", x"4B4C4C4C", x"4C4C4D4D", x"4D4D4D4D", x"4B4E4E4A", x"47474745",
									 -- x"47484847", x"47484644", x"45454443", x"44474745", x"43444547", x"46434242", x"41403F40", x"41414346",
									 -- x"44454647", x"4A4D5255", x"5658585C", x"63656568", x"6C6E7276", x"7A7D7E7E", x"7F81868B", x"8C8C8C8E",
									 -- x"8C91989B", x"9C9DA0A3", x"A1A2A6A9", x"ADB0B2B2", x"B3B5B6B7", x"BABCBBB8", x"B9BABBBC", x"BCBEC1C4",
									 -- x"C6C6C7C8", x"C9C8C9CA", x"CBCCCED1", x"D6DADDDE", x"E1E6E7E7", x"EBEDEDEF", x"EEEDEAE9", x"EAEAE9E8",
									 -- x"E6E8E9E8", x"E5E2E2E2", x"DDDDDDDC", x"DCDEDFDF", x"DDDDDDDF", x"E0DFDDDB", x"D6D7D9D9", x"D7D5D5D6",
									 -- x"D5D3D2D2", x"D3D3D4D6", x"D5D8DBDB", x"DBDDDEDF", x"E0E0DFDF", x"E0E0E0DF", x"DCDCDDDD", x"DDDBDAD9",
									 -- x"D9DDDDDB", x"DBDDD9D3", x"D0CECAC6", x"C5C5C4C2", x"C4C1BFBF", x"BEBCBBBA", x"BCBBB9B9", x"BBBCBCBB",
									 -- x"BBBBBCBE", x"BEBDBDBF", x"BABCBDBE", x"BDBCBCBC", x"BCBCBCBC", x"BDBDBDBD", x"B9B8B7B5", x"B4B4B4B4",
									 -- x"B4B1B0B2", x"B6B7B7B7", x"B8B6B3B2", x"B1AFABA8", x"A5A4A19D", x"9B9A9794", x"9594918F", x"8D8B8988",
									 -- x"8181807E", x"7D7B7A7A", x"77777675", x"7372706F", x"706E6B6A", x"69676462", x"62615F5E", x"5E5E5E5D",
									 -- x"5A5B5A58", x"57565552", x"55555350", x"4E4F4F4F", x"4C4D4D4D", x"4C4B4A4A", x"45474745", x"43444444",
									 -- x"41414141", x"403E3C3A", x"3B383536", x"37353230", x"31313030", x"302F2E2D", x"2F2E2C2A", x"2B2B2C2C",
									 -- x"2A292825", x"24262626", x"25232224", x"27282623", x"2425282B", x"2A272627", x"26292B2A", x"26242425",
									 -- x"23252221", x"24252324", x"24242423", x"23222221", x"22242422", x"21212120", x"1E1E1E1F", x"20212020",
									 -- x"20212324", x"24242525", x"282A292A", x"2D2B292C", x"2E2D2D30", x"31302F30", x"3534312F", x"2E2E2E2F",
									 -- x"2C2D2E2E", x"2D2D2E2F", x"2A2C2C2A", x"2A2E2F2D", x"2A2C2D2D", x"2B2B2C2E", x"2E2C2B29", x"2A2D3031",
									 -- x"2F2E2E2F", x"2E2D3033", x"31333332", x"31333434", x"34363736", x"36383938", x"393B3D3B", x"3737393C",
									 -- x"3B3D3F3F", x"3E3D3E3F", x"3C3D3E40", x"42434342", x"42414142", x"43444341", x"4342413F", x"41434342",
									 -- x"43434241", x"41424342", x"43434343", x"42414141", x"41414243", x"45454545", x"42454744", x"41414142",
									 -- x"4F4F4D4D", x"4E515250", x"4E4E4F50", x"51525252", x"52504F4E", x"4D4F5051", x"4C50514E", x"4C4B4B4B",
									 -- x"4C4D4C4B", x"4B4C4B49", x"494A4948", x"48494847", x"48484746", x"45454648", x"41414447", x"4949494A",
									 -- x"4A4A494B", x"4E515455", x"5757575C", x"62626369", x"71737679", x"7D7F8081", x"7F7F8185", x"888A8D90",
									 -- x"8C91979B", x"9D9EA0A2", x"A4A6A8AB", x"AEB1B5B8", x"B2B6BABB", x"BCBDBDBC", x"C0C0C0C0", x"BFC1C3C6",
									 -- x"C5C5C6C7", x"C7C7C8CA", x"CCCDCFD2", x"D6D9DCDD", x"E2E7E7E5", x"E9EDEDEF", x"EFEDECEC", x"EDEDEDEC",
									 -- x"EFEFEFED", x"EAE7E3E2", x"DFDEDCDA", x"DADBDCDC", x"DAD9D8D8", x"D8D7D5D3", x"D4D4D4D2", x"D0D0D1D2",
									 -- x"D1CFCFD0", x"D0D0D2D4", x"D6D6D7D6", x"D8DBDFE1", x"E0E0DFDF", x"E0E0DEDC", x"DDDCDCDB", x"DBDAD8D7",
									 -- x"D7D9DADA", x"D9D9D5D1", x"CFCDCAC8", x"C7C7C6C5", x"C5C1BEBF", x"BEBAB8B9", x"BAB7B5B6", x"B8B8B7B5",
									 -- x"B5B6B7B8", x"B8B8B8B9", x"B7B7B8B8", x"B9B8B7B6", x"B5B5B5B6", x"B6B7B7B7", x"B5B4B2B0", x"B0B1B1B1",
									 -- x"B1AFAEAF", x"B1B3B4B4", x"B4B2B0AF", x"AEABA7A4", x"A3A29E9A", x"98989592", x"91908D8B", x"89878584",
									 -- x"80807E7B", x"78757371", x"72727170", x"6F6D6D6C", x"6C6A6866", x"64636160", x"5D5C5B5A", x"5A5B5B5B",
									 -- x"57575552", x"51525251", x"51514F4D", x"4C4D4E4D", x"494A4A4A", x"49484747", x"43444441", x"4040403F",
									 -- x"3D3D3C3C", x"3C3C3A39", x"3A363231", x"31313131", x"33312E2D", x"2C2D2E2E", x"2C2B2B2B", x"2B2A2827",
									 -- x"25272828", x"27262423", x"24232224", x"27282725", x"24242628", x"27252425", x"27262525", x"27272523",
									 -- x"24262321", x"24242325", x"26262525", x"25242423", x"21222322", x"21212020", x"20202020", x"20202021",
									 -- x"20222425", x"25252627", x"2829292B", x"2D2C2B2E", x"2E2C2B2D", x"2F2F2E2E", x"32312F2D", x"2C2B2B2B",
									 -- x"2B2C2C29", x"2627292A", x"26282927", x"272A2C2B", x"27292A2B", x"2A2A2C2F", x"292C2D2B", x"2C2F2F2C",
									 -- x"2B2C2D2D", x"2C2C2E30", x"2F303030", x"30303131", x"34383835", x"34363736", x"37383938", x"3736383A",
									 -- x"393A3C3C", x"3C3C3C3D", x"3D3C3C3E", x"4041403E", x"3F3F3E3F", x"4040403F", x"41424140", x"3F3E3F3F",
									 -- x"4141403F", x"3F404040", x"41414141", x"41414141", x"403F3F41", x"43434342", x"43444442", x"403E3E3E",
									 -- x"53525150", x"51545452", x"52535455", x"55555555", x"55535251", x"51515253", x"4E515351", x"4F4F4F50",
									 -- x"4F4F4E4D", x"4E50504F", x"4C4E504E", x"4C4B4B4A", x"4E4D4B49", x"48494B4C", x"49494B4D", x"4D4C4B4B",
									 -- x"4F4E4D4F", x"52555554", x"595A5A5D", x"6262666E", x"75757779", x"7A7D7E80", x"7E7D7E82", x"85878A8D",
									 -- x"8E91969A", x"9D9FA0A1", x"A5A6A8A9", x"AAAEB3B8", x"B5BCC1C1", x"BFBFC0C2", x"C5C5C4C2", x"C2C3C6C8",
									 -- x"C4C6C8C9", x"CACBCCCC", x"CCCFD1D4", x"D6D8DCDE", x"E3E9EAE8", x"EBEFEFEF", x"F0EEEDEC", x"EDECEBEA",
									 -- x"EFEEEEEE", x"EFEDEAE7", x"E4E1DEDB", x"D9D9D9DA", x"D5D3D2D2", x"D2D3D2D1", x"D1D1D0CF", x"CFCECDCD",
									 -- x"CFCECECF", x"CFCECFD0", x"D5D3D2D4", x"D7DBDDDF", x"DFE0E0DF", x"E0E1DFDC", x"DEDCDAD9", x"D9D8D7D6",
									 -- x"D5D5D6D9", x"D9D5D2D1", x"CDCCCACA", x"C8C7C6C5", x"C3BFBCBD", x"BCB7B5B5", x"B6B4B2B2", x"B3B3B1AF",
									 -- x"B1B2B3B3", x"B2B2B3B3", x"B4B3B2B2", x"B3B3B2B1", x"AEAFAFAF", x"B0B0B0B0", x"AFAEABAA", x"ABACADAD",
									 -- x"AEAFAEAC", x"ACADB0B2", x"AFAFAEAD", x"ABA8A4A1", x"9E9C9995", x"9393918E", x"8C8B8886", x"84838180",
									 -- x"7E7D7B79", x"75726F6D", x"6F6F6D6C", x"6B696868", x"66656361", x"605F5E5D", x"5A585655", x"54545454",
									 -- x"51514F4C", x"4C4D4E4D", x"4D4B4947", x"494B4B48", x"46474848", x"48464443", x"3F3F3E3D", x"3E403F3C",
									 -- x"3C3B3938", x"38373736", x"3635322F", x"2D2E3031", x"33312E2C", x"2C2C2D2D", x"28282829", x"29272523",
									 -- x"23242628", x"28262322", x"22222223", x"24242424", x"26242324", x"25242324", x"26242223", x"25262524",
									 -- x"21242321", x"22212126", x"27262424", x"24242423", x"20212223", x"22212020", x"2322211F", x"1F1F2021",
									 -- x"1E212325", x"25252627", x"2927292B", x"2B2B2C2C", x"2C292729", x"2B2B2C2D", x"2E2E2E2D", x"2B292827",
									 -- x"272A2A27", x"25252626", x"23252626", x"26272828", x"25272827", x"26272A2D", x"24292A29", x"292C2B27",
									 -- x"272A2C2C", x"2B2A2C2D", x"2C2C2D2E", x"2F2E2E2E", x"30343431", x"30333534", x"34343435", x"36373635",
									 -- x"37363636", x"383A3A3A", x"3A39393A", x"3C3C3B3A", x"3D3C3B3A", x"3B3B3C3C", x"3D3F413F", x"3C393B3E",
									 -- x"3E3D3D3D", x"3D3D3D3D", x"3E3E3D3D", x"3D3D3E3E", x"3E3D3D3E", x"3F403F3E", x"43424041", x"41403E3D",
									 -- x"53555555", x"55555350", x"51525355", x"56575858", x"55555657", x"57565555", x"54565756", x"54545454",
									 -- x"53535251", x"52545554", x"4E525453", x"51505151", x"4F51504F", x"4D4D4D4C", x"4F4D4D4D", x"4D4D4D4F",
									 -- x"52515153", x"55565553", x"575A5A5B", x"5F61666F", x"76777778", x"797A7D7E", x"7E7E7F82", x"84858687",
									 -- x"8C8E9296", x"9B9D9F9F", x"A4A6A8A8", x"A9ACB2B7", x"B8BFC6C6", x"C3C2C5C7", x"C9C9C8C7", x"C6C6C9CB",
									 -- x"C7CACCCE", x"CFD1D1D1", x"CED0D3D5", x"D7D9DDE0", x"E1EAECEB", x"F0F3F1EF", x"F0EEECEC", x"EDEDECEB",
									 -- x"EEEDEDEE", x"EFEFECEA", x"E6E3DFDD", x"DAD9D9DB", x"D7D5D3D2", x"D2D2D1D1", x"CECECFD0", x"D0CECCCA",
									 -- x"CECDCECF", x"CECCCBCB", x"CFCED0D4", x"D8DAD9D9", x"DCDFDFDF", x"E0E2E1DE", x"DEDCDAD8", x"D8D7D6D5",
									 -- x"D4D2D4D9", x"D8D3D1D3", x"CDCCCCCC", x"CAC7C5C4", x"C2BFBCBB", x"BAB6B3B2", x"B3B2B1B0", x"AFAEADAC",
									 -- x"ACAEAEAD", x"ACADADAC", x"ADACABAB", x"ABABABAB", x"AAABACAC", x"ACACACAB", x"ABA9A7A7", x"A8AAAAAA",
									 -- x"ABADADAA", x"A7A8ABAD", x"AAAAA9A9", x"A7A4A09E", x"99989591", x"908F8D8A", x"87868482", x"807E7C7B",
									 -- x"77777674", x"726F6D6C", x"6C6B6A68", x"66646261", x"5F5F5E5C", x"5B595857", x"57565351", x"504F4D4C",
									 -- x"4A4B4C4B", x"4A4A4947", x"48474444", x"46494744", x"43434344", x"4443413F", x"3E3D3B3A", x"3C3D3A36",
									 -- x"3B393735", x"34333332", x"3032322F", x"2D2D2D2D", x"2F2F2E2E", x"2D2C2B2A", x"27262525", x"25252525",
									 -- x"25242526", x"26242425", x"22232323", x"23232424", x"28242223", x"24232324", x"22242524", x"21202225",
									 -- x"20232322", x"22202126", x"26242221", x"22222221", x"20202223", x"23212122", x"24221F1D", x"1E1F2020",
									 -- x"1D202223", x"22232426", x"29252729", x"27272927", x"2A282728", x"29292A2C", x"2B2B2B2B", x"29272523",
									 -- x"21262928", x"27282725", x"22232425", x"26262625", x"27282927", x"2525282A", x"25272725", x"25282827",
									 -- x"27292B2A", x"292A2A2A", x"2A2A2B2D", x"2E2D2C2C", x"2D2F302F", x"2F323333", x"35343334", x"36363532",
									 -- x"36343334", x"37393938", x"38383839", x"3A3A3A3A", x"3B3B3A39", x"39393A3B", x"3B3D3F3F", x"3B383A3E",
									 -- x"3E3D3D3E", x"3E3D3D3E", x"3F3E3C3B", x"3B3C3B3B", x"3D3D3D3E", x"3F3F403F", x"413E3D40", x"4242403F",
									 -- x"53565857", x"56565452", x"51525355", x"57595A5B", x"57585A5B", x"5B595857", x"5A5A5A5A", x"5959595A",
									 -- x"58595857", x"58595856", x"53565857", x"56575857", x"53555654", x"53535250", x"52515052", x"52535456",
									 -- x"56555556", x"57575654", x"54585757", x"5B606468", x"70727475", x"77797B7D", x"7D7D7E81", x"81828386",
									 -- x"888B8F92", x"95979A9B", x"9FA3A6A8", x"A8ABB0B5", x"B7BDC3C5", x"C6C8CBCC", x"CDCDCECD", x"CCCCCDCF",
									 -- x"CED1D4D4", x"D6D8DAD9", x"D7D7D8DA", x"DCE0E2E4", x"E3ECEDEB", x"EFF3F3F1", x"F2EFECEB", x"ECEDEDEE",
									 -- x"EDEEEEEE", x"ECEBEAEB", x"E8E4E1DF", x"DEDCDDDF", x"DDDBD9D8", x"D7D5D3D1", x"CECFD0CF", x"CDCBCACB",
									 -- x"CCCBCCCD", x"CCC9C8C8", x"CACBCED4", x"D7D6D5D6", x"D9DDDEDC", x"DCDFE0DD", x"DDDCDAD9", x"D9D8D5D2",
									 -- x"D2D2D3D4", x"D3D0CECD", x"CCCBCBCB", x"C9C5C4C4", x"C1C0BDBA", x"B8B6B3AF", x"AEAEAEAD", x"ABA9A9A9",
									 -- x"A7A9A9A8", x"A7A8A8A6", x"A6A6A6A5", x"A5A4A4A4", x"A5A6A7A8", x"A9A8A7A6", x"A8A6A4A4", x"A6A8A8A7",
									 -- x"A8AAAAA6", x"A4A5A5A4", x"A3A3A3A3", x"A19E9B99", x"9595928F", x"8E8D8A87", x"8382807E", x"7C797775",
									 -- x"7271706E", x"6D6B6968", x"67666564", x"615E5C5B", x"59595958", x"55535251", x"52514F4D", x"4C4A4947",
									 -- x"46474846", x"46464543", x"43434241", x"4243423F", x"3F3E3D3D", x"3D3D3C3B", x"3C3C3B39", x"38383633",
									 -- x"36353332", x"31313130", x"2E2F2F2D", x"2C2D2C2A", x"2C2C2C2C", x"2C2B2928", x"28262424", x"24252626",
									 -- x"27252425", x"24232425", x"23222222", x"24252524", x"24232324", x"23212022", x"1F212423", x"201E1F21",
									 -- x"21222122", x"23212025", x"24222121", x"2222201F", x"1F1F2022", x"22202022", x"211F1C1C", x"1D1F1F1E",
									 -- x"1E202222", x"21212325", x"28222528", x"24242725", x"27262728", x"28272729", x"29292827", x"26242322",
									 -- x"20242625", x"25282825", x"23222324", x"26262524", x"27282928", x"26252627", x"27262524", x"25262728",
									 -- x"28292927", x"27292A29", x"2B29292C", x"2D2C2B2C", x"2E2D2D2F", x"31313133", x"33333333", x"34343332",
									 -- x"34343435", x"36373737", x"36373838", x"3838393A", x"39393939", x"39393A3B", x"3B3B3D3E", x"3C39393B",
									 -- x"3E3C3C3E", x"3E3C3C3E", x"3E3D3C3C", x"3C3C3B3A", x"3C3D3D3D", x"3D3D3E3F", x"3E3C3C3F", x"41404040",
									 -- x"56595A59", x"58595B5B", x"58585859", x"595A5B5C", x"5B5B5B5A", x"5A595858", x"5D5B5B5B", x"5C5D5D5D",
									 -- x"5C5D5D5D", x"5C5C5A57", x"5A5A5959", x"5A5C5C5B", x"595B5C59", x"58595957", x"5858595B", x"5B5A5A5B",
									 -- x"58575757", x"58585756", x"55595755", x"5A606162", x"66696D70", x"7376797B", x"7C7B7B7C", x"7D7F8489",
									 -- x"878B8F91", x"9193969A", x"989CA2A4", x"A5A7ACB1", x"B5BAC0C4", x"C9CFD2D2", x"CFD0D2D2", x"D1D0D0D1",
									 -- x"D7DADCDC", x"DDE0E2E1", x"E4E2E0E1", x"E5E8E9E9", x"EAF0EEE9", x"EDF3F5F5", x"F8F4EEEA", x"E9EAEAEA",
									 -- x"E9ECEEED", x"EAE9EBEE", x"E9E5E2E2", x"E1E0E1E4", x"DFDEDDDD", x"DDDBD8D5", x"D2D2D0CB", x"C6C5C8CC",
									 -- x"CAC9C9CA", x"CAC8C7C8", x"CACBCED2", x"D4D3D5D8", x"D7DBDCD9", x"D8DBDCDA", x"DCDBDADB", x"DAD8D4D0",
									 -- x"CFD2D3CE", x"CCCCC9C5", x"C8C6C6C7", x"C6C2C1C3", x"BFC0BDB8", x"B5B5B1AB", x"A8AAAAA9", x"A6A4A4A5",
									 -- x"A3A5A6A4", x"A3A4A4A3", x"A1A2A3A3", x"A2A09F9F", x"9D9FA1A2", x"A3A2A1A0", x"A3A1A0A0", x"A2A4A4A3",
									 -- x"A5A7A7A4", x"A3A3A19E", x"9E9E9E9E", x"9C9A9795", x"92918F8D", x"8B8A8783", x"81807E7C", x"79767371",
									 -- x"706F6D6B", x"68666463", x"61616160", x"5E5B5958", x"57575755", x"53504E4D", x"49494848", x"47464544",
									 -- x"4444423F", x"3E40403F", x"3D3E3E3D", x"3C3C3B39", x"3D3B3838", x"38393938", x"36383938", x"36363635",
									 -- x"30303030", x"31313131", x"302F2B28", x"2A2D2C2A", x"2C2B2928", x"28292828", x"29282626", x"26262524",
									 -- x"27252526", x"25232224", x"221F1E1F", x"22242321", x"1F212425", x"221E1D1F", x"1E1E1F20", x"22211E1C",
									 -- x"1F1F1D1F", x"22201E21", x"23222122", x"2322201E", x"1E1D1E20", x"201E1F21", x"1F1C1A1A", x"1D1F1E1C",
									 -- x"20222323", x"21202225", x"26202427", x"23242825", x"22232527", x"25232224", x"27272524", x"23232323",
									 -- x"25262320", x"20252624", x"25232223", x"25262423", x"23252726", x"24232324", x"25242425", x"25252526",
									 -- x"2A2A2725", x"25292A29", x"2C2A292B", x"2C2B2B2C", x"302C2B2F", x"302E2E2F", x"2F2F2F2F", x"2E2F3032",
									 -- x"30313334", x"33323334", x"34363736", x"35343537", x"35353737", x"37373838", x"3B39383A", x"3A373534",
									 -- x"3B39393B", x"3B39383A", x"3939393A", x"3B3B3A38", x"393A3B3A", x"3938393B", x"3C3A3B3E", x"3E3C3D3F",
									 -- x"5D5A5858", x"5A5C5C5C", x"5A5B5C5C", x"5C5C5C5D", x"5B5E5D5A", x"5B60605A", x"5F5E5E5E", x"5F606060",
									 -- x"5B5C5E60", x"61605D5A", x"575A5C5D", x"5D5F6264", x"60605F5E", x"5C5A5A5A", x"5C5E6162", x"5F5C5C60",
									 -- x"5D5A595A", x"5A585758", x"5A595756", x"585B5F62", x"6564676C", x"6E6D7177", x"76777B7B", x"777A807F",
									 -- x"85888B8C", x"8F949696", x"9B9B9C9E", x"A1A5AAAD", x"B3B7BBBE", x"C3CBD0D3", x"D3D3D4D5", x"D5D5D7D8",
									 -- x"DBDEE1E5", x"E8EAEBEC", x"EDEBEAEA", x"ECEEEFEE", x"F0EFEFF0", x"F2F3F4F4", x"F5F2EEEA", x"E9E9E9E9",
									 -- x"E9EBEAE6", x"E5E7EAEB", x"EAE9E7E4", x"E3E2E1E1", x"E4E1DFE1", x"E4E4DFDA", x"D7D4D0CE", x"CCC9C9CA",
									 -- x"CACCCCC9", x"C4C3C4C7", x"CACDCFCF", x"D0D1D3D2", x"D5D6D6D5", x"D5D7D8D8", x"D8DBDDDB", x"D6D2D2D4",
									 -- x"CDCDCCCB", x"CBCAC8C7", x"C7C6C6C5", x"C4C2C0BE", x"BBBAB8B6", x"B5B2AEAB", x"A9A6A4A3", x"A3A4A3A1",
									 -- x"A0A19F9A", x"9BA0A09B", x"9B9C9C9B", x"9999999A", x"9A99999A", x"9C9C9B99", x"9E9D9A99", x"9A9DA0A1",
									 -- x"A19E9CA0", x"A3A19D9A", x"98999996", x"9493918F", x"8E8C8A89", x"8785817F", x"817E7A78", x"76736D69",
									 -- x"6B6A6866", x"64615D5B", x"5B5C5C5B", x"59565250", x"53534E4C", x"504D484B", x"47454344", x"44424142",
									 -- x"3F3D3B3A", x"393A3A3A", x"3B3A3939", x"393A3938", x"38363637", x"34353634", x"36343735", x"2E323732",
									 -- x"3030302F", x"2E2E2E2E", x"2E2B2A2C", x"2D2B2929", x"2A292928", x"27262525", x"27272624", x"26282622",
									 -- x"25262625", x"23212122", x"23212020", x"2222201E", x"22222120", x"1E1E1E1F", x"1F1E1E1E", x"1F201F1E",
									 -- x"1C1C1D1D", x"1E1F1F1F", x"23201E20", x"21202020", x"201E1D1E", x"1F1E1D1D", x"1B1A1B1C", x"1D1D1D1D",
									 -- x"1B1E2020", x"1D1D2023", x"1E212425", x"24222121", x"23232323", x"26282623", x"24242322", x"21212223",
									 -- x"25232223", x"2524221F", x"221F1F23", x"26252220", x"21212121", x"21222324", x"23222122", x"23242424",
									 -- x"25262626", x"25252526", x"27272726", x"2728292A", x"2D2B2929", x"2A2B2C2C", x"2E2D2C2D", x"2E2F2F2E",
									 -- x"2D303232", x"2F2F3236", x"33323234", x"36373737", x"34353636", x"35353637", x"37383938", x"36363739",
									 -- x"38393B3B", x"39383839", x"3B3A3939", x"3A393837", x"39393938", x"3838393A", x"3B3B3B3B", x"3A3A3C3C",
									 -- x"5D5C5B5B", x"5C5D5C5C", x"5D5D5E5F", x"5F5E5D5C", x"5E5E5E5E", x"60626260", x"5F606161", x"5F5F6162",
									 -- x"61616061", x"615F5D5B", x"5D5E6061", x"61636567", x"66646160", x"5F5E5D5C", x"61606161", x"605E6063",
									 -- x"615F5E60", x"605F5F60", x"5F5E5C5B", x"5B5D5E60", x"60626566", x"676A6D6F", x"6E707476", x"757A7F7F",
									 -- x"7E83888A", x"8C8F908F", x"96989B9D", x"A0A3A7AA", x"AFB3B8BB", x"BFC6CCCF", x"D3D4D5D6", x"D7D9DADB",
									 -- x"DDDFE2E6", x"E9ECEDED", x"EEEFF0F1", x"F2F2F1F0", x"F2F1F1F1", x"F1F2F2F3", x"F2F0EEEC", x"ECECECEC",
									 -- x"E8E8E7E4", x"E4E6E8E8", x"E9E8E7E6", x"E5E4E3E3", x"E0E1E3E3", x"E1DFDEDD", x"D9D6D3D2", x"D0CECDCE",
									 -- x"C8C9C9C8", x"C6C4C4C5", x"C6CACECF", x"CFD0D1D1", x"D2D3D4D4", x"D5D6D7D6", x"D5D7D7D6", x"D4D1D0D0",
									 -- x"CFCDCBCA", x"C9C8C7C7", x"C4C4C4C4", x"C3C0BDBB", x"B8B6B5B3", x"B2AFABA9", x"A8A6A2A1", x"A1A09F9D",
									 -- x"9D989799", x"9996979B", x"96979797", x"95949494", x"94959595", x"95949494", x"96959594", x"9596989A",
									 -- x"9B98989B", x"9D9B9896", x"91929290", x"8F8F8E8C", x"88868483", x"82807D7B", x"77757372", x"72716D6A",
									 -- x"67666463", x"615E5B59", x"55565656", x"54524F4D", x"4C4B4848", x"4A474445", x"44424141", x"403E3D3D",
									 -- x"3B3A3837", x"36373737", x"38373535", x"35363636", x"38353535", x"3130312E", x"33313433", x"2E30332F",
									 -- x"2F2F2E2D", x"2C2B2C2C", x"2C2A2A2D", x"2E2B2827", x"2A292726", x"27262524", x"24242322", x"22242320",
									 -- x"23232322", x"21212122", x"21201F1F", x"1F1F1E1D", x"2020201F", x"1E1E1E1F", x"1F1E1D1C", x"1D1E1E1D",
									 -- x"1B1C1D1E", x"1E1E1E1E", x"22201F1F", x"1F1E1E1F", x"1C1B1B1E", x"1F1D1B1A", x"1C1B1C1C", x"1D1D1D1C",
									 -- x"1B1D1E1D", x"1C1B1D20", x"1E202123", x"23232323", x"24242222", x"24262624", x"22232322", x"21212122",
									 -- x"24232222", x"22222120", x"221F1F22", x"24242120", x"20201F1F", x"20202122", x"22212122", x"24242423",
									 -- x"24242525", x"24242525", x"24252626", x"2526282B", x"2B2A292A", x"2C2D2D2D", x"2D2C2C2C", x"2D2E2E2D",
									 -- x"2B2D2E2F", x"2F2F2F30", x"31303031", x"32333232", x"35353535", x"35353535", x"35343435", x"35353534",
									 -- x"34363737", x"36353738", x"39383838", x"3A3B3B3A", x"38383837", x"36353637", x"36373838", x"3839393A",
									 -- x"5E5F6060", x"5F5E5E5D", x"61626263", x"6362615F", x"66636265", x"66646364", x"60636665", x"62616467",
									 -- x"68666462", x"6261605F", x"60616162", x"64656667", x"6A676361", x"6262605E", x"65636262", x"63636465",
									 -- x"64636364", x"64646464", x"63636261", x"605F5F5F", x"5D636562", x"62676967", x"66696D6F", x"72777A7A",
									 -- x"797E8486", x"87898B8C", x"8F93989B", x"9C9FA3A6", x"AAAEB2B5", x"BAC0C6C9", x"CECED0D2", x"D5D7D9D9",
									 -- x"DBDDE0E5", x"EAEEF0F0", x"F0F1F3F3", x"F3F2F1F0", x"F0F0F0EE", x"ECEBEBEC", x"E9E9E9E9", x"EAEBEAEA",
									 -- x"E5E5E4E2", x"E3E4E5E4", x"E6E7E7E7", x"E6E5E4E3", x"DFE1E3E4", x"E3E2E1E1", x"DBD8D6D6", x"D4D1D0D0",
									 -- x"CAC8C6C4", x"C4C3C3C2", x"C6CBCFD0", x"CFCECDCC", x"CDD0D1D1", x"D1D3D2D0", x"D4D4D4D4", x"D4D2D0CE",
									 -- x"D0CECAC7", x"C6C6C6C6", x"C2C2C3C3", x"C2BEBAB7", x"B5B4B3B3", x"B2AFABA8", x"A7A4A19F", x"9F9E9C9A",
									 -- x"97949395", x"938F9095", x"90919291", x"908F8F8F", x"8D8F9090", x"8E8C8C8D", x"8E8F9090", x"8F909193",
									 -- x"94939395", x"95949393", x"8F908F8C", x"8A8A8886", x"8382807E", x"7E7C7977", x"71706F6E", x"6D6B6867",
									 -- x"62605F5D", x"5C5A5857", x"4F4F4F4F", x"4E4C4B4A", x"48444445", x"4342413F", x"3F3E3D3D", x"3B393737",
									 -- x"37363534", x"34343433", x"35343231", x"32323333", x"38353534", x"302F2F2C", x"2F2D3031", x"2F31322D",
									 -- x"2F2E2E2D", x"2D2D2D2D", x"2C2A2A2B", x"2C2A2827", x"2A272525", x"26272523", x"24252422", x"22232322",
									 -- x"24232221", x"21212222", x"20201F1F", x"1E1E1D1D", x"1E1F1F1E", x"1D1D1D1E", x"1F1D1B1A", x"1B1B1C1C",
									 -- x"1B1C1D1E", x"1E1E1D1D", x"201F1E1F", x"1E1C1C1E", x"1B19191B", x"1C1B1918", x"1B1B1B1B", x"1C1C1B1A",
									 -- x"1A1B1C1C", x"1C1C1D1E", x"1F1F1E1F", x"21222323", x"23232222", x"23252422", x"21212222", x"21212121",
									 -- x"22222221", x"1F1F2021", x"211F1F21", x"22212021", x"21212020", x"20212122", x"21212222", x"23232221",
									 -- x"22222323", x"23232425", x"23252626", x"2424272A", x"2828292A", x"2B2C2B2A", x"2C2B2B2B", x"2C2D2D2C",
									 -- x"2C2B2C2D", x"2F302E2C", x"31302F2F", x"30302F2F", x"35333231", x"32333232", x"34323133", x"36373431",
									 -- x"30323233", x"33343638", x"39383736", x"37383838", x"36363635", x"34333333", x"34353739", x"39393939",
									 -- x"60626565", x"63616162", x"66676868", x"67656565", x"69686769", x"6A6A6868", x"64676867", x"6564676A",
									 -- x"6A696765", x"64646464", x"63626263", x"65676767", x"68676462", x"6262615F", x"62636465", x"66666565",
									 -- x"66656566", x"66666665", x"66666564", x"63626262", x"60646664", x"63666664", x"65696A6B", x"6F717171",
									 -- x"767A7E80", x"8083888B", x"8B8F9396", x"97999FA3", x"A5A8ACB0", x"B5BBC1C4", x"C5C7C8CA", x"CED2D3D2",
									 -- x"D5D7DAE0", x"E8EEF1F1", x"F1F1F1EF", x"EDECEDEE", x"EBECECE9", x"E5E3E4E5", x"E3E2E3E4", x"E5E6E5E5",
									 -- x"E2E1E0E0", x"E1E3E3E1", x"E2E3E5E6", x"E6E5E4E3", x"E2E0DFE1", x"E4E6E4E1", x"DCD9D7D7", x"D5D2CFCE",
									 -- x"CECAC5C1", x"C0C0C0C0", x"C6C9CCCD", x"CECFCDCA", x"CDCFD0CF", x"CFD0CFCD", x"D4D4D5D5", x"D5D3D2D1",
									 -- x"D0CDCAC7", x"C5C5C5C4", x"C3C3C3C2", x"C0BCB8B5", x"B6B6B7B8", x"B7B4AFAB", x"A7A4A1A0", x"A09F9C9A",
									 -- x"94979692", x"90918F8A", x"8B8B8B8A", x"8A898A8A", x"8A8B8B8B", x"89888888", x"87888A8A", x"89888A8C",
									 -- x"8C8C8D8E", x"8D8B8C8E", x"8C8D8B88", x"86858381", x"7F7D7B7A", x"79777573", x"6E6E6D6B", x"68656463",
									 -- x"5D5C5A58", x"57555453", x"4D4C4B4A", x"49484747", x"48414345", x"3F3E3F3A", x"39393939", x"37353333",
									 -- x"34343332", x"32323231", x"32323131", x"31313131", x"34323333", x"2F2F2F2C", x"2D2C2D30", x"31333230",
									 -- x"2F2E2E2E", x"2F2F2F2F", x"2E2C2928", x"28282828", x"27262424", x"24252524", x"25252523", x"22232424",
									 -- x"25232121", x"2121201F", x"20212120", x"1F1E1E1E", x"1E1E1E1D", x"1C1B1B1C", x"1D1C1B1B", x"1A1B1B1B",
									 -- x"1C1C1C1D", x"1D1D1D1D", x"1C1C1D1E", x"1D1B1D1F", x"1E1B1818", x"19181819", x"19191919", x"1A1A1919",
									 -- x"1B1B1B1C", x"1D1E1F1F", x"201E1D1E", x"20212121", x"21222323", x"2424221E", x"20212020", x"1F1F2021",
									 -- x"2020201F", x"1E1E1E1F", x"1F1E1F20", x"1F1E1F21", x"21212020", x"20202121", x"20202021", x"21212020",
									 -- x"20212222", x"22222324", x"25262625", x"25252627", x"26262728", x"28282727", x"292A2A2A", x"2B2B2B2B",
									 -- x"2C2B2A2C", x"2E2E2C2A", x"2F2F2F2E", x"2E2E2D2D", x"32302D2E", x"2F30302E", x"32302F31", x"34353331",
									 -- x"2F303030", x"31333638", x"39383635", x"35353637", x"35363635", x"34333333", x"3435383A", x"3A393938",
									 -- x"63656767", x"65656668", x"686B6C6B", x"6867696C", x"686B6C6B", x"6D71716D", x"6B6A6969", x"68676767",
									 -- x"6A696867", x"66656565", x"66666566", x"68696969", x"64676865", x"63636362", x"61646666", x"66666768",
									 -- x"68686869", x"6A6B6A69", x"69686665", x"64646565", x"65656666", x"66656464", x"656A6A69", x"6D6E6B6D",
									 -- x"7074787A", x"7B7D8287", x"878A8E8F", x"90949AA0", x"A0A3A7AC", x"B0B6BBC0", x"BFC1C3C4", x"C8CCCDCB",
									 -- x"D0D1D5DB", x"E3EAEEF0", x"EEEFEEEC", x"E9E8E8E9", x"E7E8E8E5", x"E1DFDFE0", x"E1E0DFDF", x"E0E1E1E0",
									 -- x"DDDCDCDD", x"DFE0E0DF", x"DFE0E2E4", x"E5E5E4E3", x"E1DEDCDD", x"E0E2E1E0", x"DDDAD7D7", x"D5D1CDCC",
									 -- x"CDCBC8C4", x"C2C1C0C0", x"C0C1C2C5", x"CACECECB", x"CDCECECD", x"CECFCFCD", x"D2D3D5D4", x"D3D2D2D3",
									 -- x"D0CECCC9", x"C8C7C6C5", x"C6C5C3C0", x"BDBAB7B4", x"B8B9BBBD", x"BDB9B2AE", x"A8A6A2A1", x"A09F9C99",
									 -- x"95979592", x"92938E86", x"87868584", x"84848585", x"86868585", x"86858482", x"81808182", x"817F8084",
									 -- x"84848586", x"84828386", x"83848381", x"8080807E", x"7A787573", x"72716E6C", x"69696966", x"63616060",
									 -- x"5A595654", x"5351504E", x"4B4A4846", x"45434242", x"453F4041", x"3C3A3B37", x"34363636", x"34333231",
									 -- x"31302F2F", x"2F302F2F", x"30303132", x"3231302F", x"302E3030", x"2D2D2E2B", x"2E2D2D2E", x"31313031",
									 -- x"302F2E2E", x"2E2E2E2D", x"2C2C2A28", x"27262524", x"23242424", x"22222425", x"23222221", x"20202123",
									 -- x"21201F1F", x"201F1D1B", x"20202020", x"1F1E1F1F", x"1C1D1D1D", x"1C1B1B1C", x"1B1B1C1C", x"1C1B1B1B",
									 -- x"1C1C1B1B", x"1B1C1D1D", x"1B1C1D1E", x"1D1C1D1F", x"201C1919", x"19181819", x"19181819", x"1A1A1A19",
									 -- x"1D1C1B1C", x"1E1F1F1F", x"1F1E1E1F", x"21222120", x"21222221", x"2122211E", x"21201F1E", x"1D1E2021",
									 -- x"1F1E1E1E", x"1E1E1D1C", x"1E1D1E1E", x"1E1C1D20", x"1F1E1E1D", x"1D1E1E1F", x"201F1F1E", x"1D1E1F1F",
									 -- x"20202122", x"22222323", x"26242223", x"25262423", x"24242425", x"25252626", x"27272828", x"28282828",
									 -- x"28282828", x"28282929", x"2B2C2C2B", x"2B2B2B2B", x"2F2D2B2C", x"2E2F2E2D", x"2E2D2D2D", x"2D2E3030",
									 -- x"31303030", x"30313233", x"34343333", x"34353839", x"35363636", x"35353535", x"33353739", x"38373636",
									 -- x"65676969", x"68686A6C", x"6B6D6E6D", x"6A6A6D71", x"6E72726F", x"7075746E", x"726F6C6A", x"6B6A6764",
									 -- x"696A6A69", x"67666666", x"69696969", x"696A6A6A", x"656A6D6A", x"67676766", x"66686866", x"66686B6D",
									 -- x"696A6B6B", x"6C6E6E6C", x"6C6B6967", x"66666767", x"68676667", x"67656465", x"646C6A68", x"6E6D6A6E",
									 -- x"6C70757A", x"7B7C7F83", x"83868889", x"8B8F959A", x"9C9EA1A6", x"AAAFB4B9", x"B7BBBEBE", x"C0C4C6C4",
									 -- x"CBCDD1D6", x"DCE2E7EA", x"E9EBECEC", x"EAE7E5E3", x"E2E2E3E1", x"DEDBDADA", x"DDDCDADA", x"DADADADA",
									 -- x"D9D7D7D9", x"DADADBDC", x"DCDDDFE1", x"E2E3E3E3", x"DFE0E0DE", x"DBDBDEE1", x"DEDAD6D5", x"D5D1CECD",
									 -- x"CBCBCBCB", x"C9C7C5C3", x"C1C0BEBF", x"C3C7C7C4", x"C5C7C8C8", x"C9CCCCCC", x"CDCED0CF", x"CECED0D2",
									 -- x"D2D1CECC", x"CBC9C7C6", x"C7C5C2BE", x"BCB9B7B5", x"B9BABCBE", x"BEBAB3AF", x"AAA8A4A1", x"A09D9A97",
									 -- x"97919094", x"96908A89", x"87868483", x"83838383", x"817F7E7F", x"807F7D7B", x"7D7A7879", x"7977787A",
									 -- x"7C7D7E7F", x"7D7C7D80", x"7D7E7D7A", x"79797977", x"7573706E", x"6D6B6967", x"66656360", x"5D5A5858",
									 -- x"57555351", x"4F4D4B4A", x"48464442", x"403F3E3E", x"3D3A3A3A", x"37353535", x"30333432", x"31313130",
									 -- x"2F2E2D2D", x"2D2E2E2E", x"2F313333", x"33313030", x"32303131", x"2E2E2E2C", x"2F302D2C", x"302E2C30",
									 -- x"33322F2E", x"2E2E2C2B", x"282A2A29", x"27262320", x"21232524", x"21202223", x"22202020", x"201F2021",
									 -- x"1D1E1F20", x"201F1D1C", x"1E1E1E1E", x"1E1E1E1E", x"1B1C1C1D", x"1C1C1C1D", x"1A1B1D1D", x"1D1C1B1B",
									 -- x"1C1B1B1A", x"1B1C1C1D", x"1C1C1D1E", x"1D1B1C1D", x"1E1B1B1C", x"1D1A1716", x"1A1A1A1A", x"1B1C1B1A",
									 -- x"1D1D1C1C", x"1D1D1D1D", x"1E1E1F20", x"21222221", x"2222201E", x"1D1F2120", x"20201E1D", x"1C1C1E20",
									 -- x"1D1D1D1D", x"1E1E1C1A", x"1D1C1C1D", x"1D1B1C1E", x"1E1D1D1D", x"1D1D1E1E", x"1F1F1E1C", x"1C1C1E20",
									 -- x"1F202121", x"21212122", x"221F1D1F", x"23252320", x"22222323", x"23242628", x"24252627", x"26262626",
									 -- x"26272827", x"26262729", x"29292A2A", x"2A2A2A2B", x"2C2B2A2B", x"2D2D2C2B", x"2B2C2C2B", x"292A2D30",
									 -- x"3130302F", x"2E2E2D2D", x"3130302F", x"2F313335", x"35353636", x"36363637", x"35373838", x"38373636",
									 -- x"67686A6B", x"6B6B6D6E", x"6E6F6F70", x"70717374", x"76777776", x"76777571", x"7773706F", x"706F6C69",
									 -- x"6A6B6C6C", x"6B6A6B6B", x"6D6D6E6C", x"6B6A6B6C", x"6B6F706D", x"6B6C6C6A", x"6D6E6C6A", x"6A6C6E6E",
									 -- x"6B6D6D6D", x"6E6F6E6C", x"6E6D6B6A", x"696A6A6A", x"6A6C6B68", x"68696966", x"656F6C69", x"6E6D6970",
									 -- x"6E6F7478", x"7A7B7D80", x"7E808486", x"898C8F92", x"98999CA1", x"A4A7ABB0", x"B0B6BAB9", x"B9BDBFBF",
									 -- x"C5C8CCD0", x"D5DAE0E5", x"E5E5E7E8", x"E7E6E3E1", x"DEDFDFDF", x"DDDAD8D6", x"D7D6D5D4", x"D4D4D4D3",
									 -- x"D4D3D3D4", x"D4D3D5D7", x"D9D9DADB", x"DDDFE0E1", x"DEE0E1DF", x"DCDBDDDF", x"DCD7D4D3", x"D4D2D1D0",
									 -- x"CFCECDCE", x"D0CFCCC9", x"C8C7C4C0", x"BFC0C0BE", x"BEC1C3C4", x"C6C8C9C7", x"CACACACA", x"CCCECFD1",
									 -- x"D4D2CFCD", x"CBC9C7C6", x"C4C2BFBD", x"BAB8B6B5", x"B8B9BABB", x"BBB7B2AE", x"ACA9A5A3", x"A19E9A96",
									 -- x"97918F92", x"938E8989", x"87858483", x"82817F7E", x"7A7A7979", x"78777675", x"77727072", x"72706F70",
									 -- x"72737576", x"76757679", x"77777673", x"7171716F", x"6F6D6A69", x"68666563", x"61605D5A", x"57545251",
									 -- x"52514F4E", x"4C4A4745", x"4342413F", x"3E3D3C3C", x"39383533", x"33302F32", x"2D30312F", x"2D2E2F2F",
									 -- x"32312F2F", x"2F303131", x"31333536", x"35343333", x"36333333", x"2F2F302D", x"2E312D2D", x"302D2A30",
									 -- x"34312F2E", x"2E2E2C2A", x"26282927", x"25252321", x"22232423", x"21201F1F", x"23201F21", x"22212020",
									 -- x"1D1E1F20", x"1F1E1D1D", x"1D1C1C1D", x"1E1F1F1E", x"1C1D1E1E", x"1D1C1C1C", x"1B1C1D1D", x"1C1B1B1C",
									 -- x"191A1A1B", x"1C1C1C1C", x"1C1B1B1D", x"1D1C1B1C", x"1C1A1A1C", x"1D1A1817", x"1B1B1B1B", x"1C1C1B1A",
									 -- x"1C1C1C1C", x"1C1D1D1E", x"1C1D1E1E", x"1E1E1F20", x"2021201E", x"1D1F201F", x"1F1F1E1D", x"1C1C1C1D",
									 -- x"1C1D1D1D", x"1C1B1B1C", x"1C1B1B1C", x"1C1B1B1C", x"1D1D1C1C", x"1D1D1E1F", x"1E1E1E1D", x"1C1D1E20",
									 -- x"1E1F2020", x"1F1F2020", x"1F1D1C1E", x"22242220", x"20212222", x"22232526", x"21232525", x"24242424",
									 -- x"24262727", x"26252728", x"26272828", x"2828292A", x"28292A2A", x"2A2A2929", x"292A2A29", x"28282B2D",
									 -- x"2E2E2E2F", x"2F2E2D2B", x"2F2F2F2E", x"2D2D2F30", x"34343434", x"34343536", x"36373737", x"36353636",
									 -- x"68696B6D", x"6D6D6D6D", x"72717173", x"77787876", x"7675767A", x"7C7B7A7A", x"78767473", x"74757371",
									 -- x"6B6D6E6F", x"6F707172", x"72737472", x"6F6D6E6F", x"7072716D", x"6D6F6F6B", x"7171706E", x"7072706C",
									 -- x"70727270", x"70706E6B", x"6D6D6D6C", x"6C6D6D6D", x"6D72706A", x"696F6F69", x"68726F6A", x"6E6B686F",
									 -- x"706F7073", x"76777A7E", x"797D8185", x"888A8B8C", x"9696999D", x"9FA1A5AA", x"ADB4B9B8", x"B7BBBEBE",
									 -- x"BEC2C7CB", x"CFD5DCE1", x"E2E1E0E1", x"E2E3E2E1", x"E0E0E0E0", x"DFDCD9D6", x"D3D3D2D2", x"D2D2D1D1",
									 -- x"D2D1D1D1", x"D0CED0D3", x"D5D5D6D7", x"D8DBDDDE", x"DDDCDBDC", x"DEDEDDDB", x"DAD5D1D1", x"D3D3D2D2",
									 -- x"D6D1CDCE", x"D2D4D2CE", x"CCCDCAC5", x"C0BFC0C0", x"BDC0C3C5", x"C6C8C8C6", x"C9C8C6C8", x"CCD0D1D1",
									 -- x"D4D2CECB", x"C9C7C5C4", x"C1C0BDBB", x"BAB8B6B5", x"B9B8B8B8", x"B7B5B1AE", x"ACA9A6A4", x"A29F9C98",
									 -- x"9496938D", x"8C8E8C86", x"84828181", x"7F7D7A77", x"76777876", x"73717171", x"706A686A", x"6C686666",
									 -- x"68686B6D", x"6E6D6F71", x"6D6D6C6B", x"6A6C6C6B", x"69676463", x"6261605E", x"5A595755", x"55545352",
									 -- x"4E4E4C4B", x"4A474543", x"40403F3E", x"3D3C3C3C", x"383A3431", x"322E2B31", x"2C2F302D", x"2B2C2D2D",
									 -- x"37353433", x"33343536", x"35363838", x"37363636", x"36333332", x"2E2E2F2D", x"2C302E2E", x"322E2B33",
									 -- x"2F2D2B2B", x"2C2C2A29", x"28282622", x"21232524", x"24242323", x"22201D1C", x"221F1E20", x"22211F1F",
									 -- x"1D1E1F1E", x"1C1A1B1B", x"1E1C1B1D", x"1F21201E", x"1F1F1F1F", x"1D1B1A1A", x"1C1D1D1C", x"1B1A1B1C",
									 -- x"17191B1C", x"1D1D1C1B", x"1B19191C", x"1E1D1C1C", x"1C191819", x"1A191919", x"1B1B1B1B", x"1B1B1A19",
									 -- x"1A1B1C1D", x"1D1E1F21", x"1B1C1D1C", x"1A1A1B1C", x"1C1F2121", x"20201E1C", x"1E1E1F1E", x"1D1C1B1B",
									 -- x"1B1D1E1C", x"1A191B1E", x"1C1A1A1C", x"1C1B1A1B", x"1A1A1A1A", x"1B1C1D1D", x"1D1E1F1E", x"1D1D1F20",
									 -- x"1E1E1F1F", x"1E1E1E1F", x"1F1E1E1F", x"21222120", x"1F202121", x"20202223", x"20222424", x"23222323",
									 -- x"21222324", x"24242424", x"23242525", x"25252627", x"26272829", x"28262625", x"25262726", x"26262728",
									 -- x"2A2B2D2F", x"31302F2E", x"2E2F2F2F", x"2F303335", x"33333332", x"32323435", x"34343433", x"32323334",
									 -- x"6C6B7170", x"70726F71", x"73717377", x"7776777B", x"76787A7B", x"7D7F8081", x"79787A7C", x"7C777372",
									 -- x"71747473", x"74777570", x"72747778", x"76737376", x"74737172", x"74757473", x"72767672", x"71747470",
									 -- x"7372706F", x"6F6F7070", x"6E6C6D6F", x"6E6A6A6D", x"6B6F706E", x"71767570", x"7274726D", x"696C7072",
									 -- x"70707070", x"73797C7C", x"7C7C7E80", x"84888A8A", x"8E919497", x"9A9EA3A6", x"AAA8AAB0", x"B4B6B7B9",
									 -- x"C0BFC1C7", x"CDD1D5D9", x"DFDEDDDD", x"DEDFDFDF", x"E0DEDDDD", x"DDDCD8D5", x"D2D3D0CB", x"CACDCECB",
									 -- x"CBCBCCCD", x"CCCBCCCF", x"CDCED0D1", x"D2D5D7D9", x"D6D7D8D9", x"D9D9D8D8", x"D8D7D5D4", x"D3D4D5D5",
									 -- x"D2D3D1CF", x"D1D7D7D4", x"D0CECAC4", x"C1C1C2C1", x"C1C3C4C4", x"C7C9C9C6", x"CCCCC8CC", x"D1D1D5D1",
									 -- x"D1CECBC8", x"C8C8C7C6", x"C6C0BBBA", x"BAB7B4B2", x"AEB1B4B5", x"B3B0AEAD", x"A5A5A2A0", x"A09F9A94",
									 -- x"94928E8B", x"8B8C8986", x"8381807F", x"7D787575", x"73717070", x"6F6C6867", x"69676563", x"62616060",
									 -- x"60616365", x"67686765", x"66656363", x"63626365", x"64625F5B", x"5B5B5955", x"56565451", x"4F4F4E4D",
									 -- x"4D494646", x"45444343", x"403D3C3D", x"3B383636", x"3B363332", x"312F2E2E", x"2E2E2F31", x"31303132",
									 -- x"38383635", x"383B3A36", x"3C3E3E3D", x"3C3B3937", x"38363432", x"302E2D2D", x"312F2F30", x"3232312E",
									 -- x"2E2E2D2A", x"2A2C2B28", x"2A272423", x"24252525", x"23232324", x"2524211F", x"231F1E21", x"22201E1F",
									 -- x"1C1C1A18", x"1A1E1E1B", x"181B1B19", x"1A1C1C19", x"1C1D1D1C", x"1B1B1C1D", x"1F1B181A", x"1C1D1C1D",
									 -- x"1C1D1C19", x"191A1A17", x"1E19181B", x"1D1B1A1B", x"181F1E18", x"171D1F1B", x"171A1B1A", x"191A1B1B",
									 -- x"1C1E201F", x"1E1C1C1C", x"1D1D1C1D", x"1F1E1D1B", x"1B1E201F", x"1C1A1C1E", x"1F1E1E1E", x"1F1F1E1D",
									 -- x"1A1B1C1B", x"1A19191A", x"191C1C1A", x"19191918", x"19191A1C", x"1C1A1A1B", x"1E1E1D1D", x"1D1D1D1D",
									 -- x"1D1D1E1E", x"1E1D1E1F", x"1B1E1E1C", x"1E21201B", x"2021201E", x"1E212120", x"201F1E1E", x"20232422",
									 -- x"1F202123", x"23242525", x"24232221", x"22242627", x"23232427", x"26252629", x"2A272425", x"28292725",
									 -- x"28292A2A", x"29292A2B", x"282A2D2D", x"2C2C2F32", x"3233322E", x"2E31322F", x"31343433", x"33303239",
									 -- x"6B6A6F6E", x"6E706D6F", x"70707276", x"78787877", x"75797D7D", x"7C7B7B7C", x"7C7B7C7E", x"7D797676",
									 -- x"72737576", x"78797875", x"7576787A", x"7A797B7E", x"7A797879", x"7B7C7B79", x"7B7B7975", x"75787875",
									 -- x"72717171", x"72737374", x"73717172", x"72706F6E", x"6F707071", x"73747473", x"73747471", x"6F727475",
									 -- x"73747575", x"787E8183", x"7D7E7F81", x"83868889", x"8B8D9092", x"94979C9F", x"A5A4A6AB", x"B0B2B3B5",
									 -- x"BBBBBDC3", x"C8CCCFD2", x"D9D8D8D8", x"D8D8D8D9", x"D9D9D9D9", x"D9D7D6D5", x"CFD0CDC8", x"C7CACAC7",
									 -- x"C8C7C7C8", x"C9C8C9CA", x"CACCCFD1", x"D2D2D3D3", x"D3D3D3D3", x"D3D3D4D4", x"D4D4D3D2", x"D2D2D3D4",
									 -- x"D1D2D1CF", x"D2D7D8D5", x"D1CFCBC5", x"C2C3C3C2", x"C5C5C4C3", x"C5C8C9C7", x"C9CBC9CD", x"CECDD0CD",
									 -- x"CAC9C7C7", x"C8C8C7C6", x"C4BFBAB9", x"B9B7B5B4", x"B0B1B3B3", x"B1AEABAA", x"A09F9D9A", x"9A999692",
									 -- x"908E8A88", x"88898683", x"817E7C7A", x"77737171", x"6E6C6A6B", x"6A676564", x"64626160", x"605F5F5E",
									 -- x"605F5D5D", x"5D5F5F5F", x"5E5D5C5C", x"5B5A5C5F", x"5E5E5C58", x"57575451", x"53524F4C", x"4B4C4B49",
									 -- x"47454444", x"43424244", x"3D3B393A", x"3A373433", x"36333131", x"32323234", x"312F2E30", x"31333437",
									 -- x"393C3D3C", x"3B3E4143", x"44444443", x"42413D39", x"34333130", x"2F2F2E2D", x"30303031", x"33343332",
									 -- x"2A2F332F", x"2B2A2C2D", x"26262727", x"26242322", x"23222222", x"22221F1E", x"21222221", x"1F1F1F1F",
									 -- x"1D1D1B1A", x"1C1E1D1A", x"1B1C1C1B", x"1B1C1B1A", x"1B1C1D1D", x"1D1C1C1C", x"1D1A181A", x"1C1B1A19",
									 -- x"1A1B1A19", x"191A1917", x"201B1514", x"15171B1D", x"191D1D18", x"171B1C1A", x"191B1C1A", x"1A1C1C1C",
									 -- x"1C1C1C1C", x"1B1A1A1A", x"1D1C1B1C", x"1D1D1C1B", x"1A1C1E1D", x"1C1B1C1E", x"1E1D1C1C", x"1D1D1D1C",
									 -- x"1A1B1B1B", x"1A19191A", x"1B1B1A19", x"1A1C1C1A", x"1918191B", x"1B1A1A1B", x"1D1D1D1D", x"1D1D1D1C",
									 -- x"1E1E1E1E", x"1D1D1C1C", x"1D1F1F1D", x"1E21201D", x"1D1F1F1E", x"1E1F1F1E", x"1F201F1E", x"1F212120",
									 -- x"1F1F1F20", x"21212121", x"21202020", x"20222324", x"24232324", x"23232528", x"27252324", x"25262523",
									 -- x"27282A2A", x"29292A2B", x"2A2B2B2B", x"2B2C2D2E", x"2E303130", x"2E2E3030", x"32353534", x"34313137",
									 -- x"6C6B6F6D", x"6D6F6C6F", x"70706F71", x"74777673", x"72777B7C", x"79767677", x"77777879", x"78767474",
									 -- x"7676777A", x"7B7A7877", x"7C7B7B7C", x"7C7B7D80", x"7F7E7E7F", x"8181807F", x"8583807F", x"7F7E7D7B",
									 -- x"7A797979", x"79797978", x"77777575", x"76777571", x"73727273", x"73717275", x"77787777", x"787A7A79",
									 -- x"797B7C7B", x"7B7E8182", x"80808182", x"83848688", x"8A8C8E90", x"9194989B", x"9E9EA0A5", x"A9ABADAF",
									 -- x"B5B5B8BE", x"C2C5C7C8", x"CCCECFD0", x"D0D0D2D4", x"D0D1D2D2", x"D1D1D1D2", x"CCCCC9C5", x"C4C6C5C3",
									 -- x"C6C4C2C5", x"C7C6C6C6", x"C7C9CBCC", x"CDCCCCCC", x"D1D0CFCE", x"CECFCFD0", x"CFCFCECE", x"CECECECE",
									 -- x"CECFCECE", x"D0D5D6D4", x"D2D1CDC8", x"C5C4C4C3", x"C4C4C3C3", x"C4C7C8C7", x"C6CAC9CC", x"CBC8CBC8",
									 -- x"C5C5C6C8", x"CACBCAC9", x"C9C4BFBD", x"BBB8B5B4", x"B2B1B0AE", x"ADAAA7A5", x"9E9D9B98", x"96959390",
									 -- x"8D8C8986", x"86868480", x"7D7A7774", x"726F6D6D", x"68666465", x"64626160", x"5E5D5B5A", x"5A5A5959",
									 -- x"5A585554", x"54555657", x"55545556", x"5555575A", x"58595957", x"5654514F", x"52504C4A", x"4A4C4A47",
									 -- x"45454545", x"43414245", x"3E3C3B3B", x"3B383634", x"38363433", x"33333334", x"35323031", x"3335383B",
									 -- x"3B3E403F", x"4043484A", x"4B4B4A49", x"4948433D", x"35353331", x"32343330", x"32333436", x"37383837",
									 -- x"3333312F", x"2E2E2D2B", x"26282A29", x"27242222", x"24232221", x"21201F1E", x"2025251F", x"1B1D1F1F",
									 -- x"1E1E1D1D", x"1D1E1D1A", x"1D1B1B1C", x"1C1B1B1C", x"1A1B1C1D", x"1E1E1C1A", x"1D1B1A1D", x"1E1D1A19",
									 -- x"191A1A19", x"19191816", x"1B1B1917", x"181A1A19", x"181A1B19", x"17181919", x"191A1A1A", x"1B1C1C1B",
									 -- x"1D1C1B1A", x"1A1A1A1A", x"1C1A1919", x"1B1B1B1A", x"1A1B1B1B", x"1B1B1C1D", x"1D1C1B1B", x"1C1D1D1D",
									 -- x"1A1B1B1A", x"1A19191A", x"1D1B1918", x"1A1D1D1A", x"1A181719", x"1B1B1A1A", x"1B1B1C1C", x"1C1C1C1B",
									 -- x"1D1D1C1D", x"1D1D1B19", x"1B1D1D1B", x"1B1D1E1D", x"1A1C1D1C", x"1C1D1D1B", x"1E1F1F1E", x"1D1E1E1D",
									 -- x"1F1E1D1E", x"1F1F1E1D", x"1F1F1F20", x"20212122", x"22222223", x"23222324", x"25242323", x"24242423",
									 -- x"26272828", x"2828292B", x"2D2B2929", x"2A2B2B2A", x"2A2D2F30", x"2E2B2D31", x"30323232", x"34312F33",
									 -- x"6F6D716E", x"6E706D70", x"71716E6A", x"6C717370", x"70727576", x"75737273", x"76777879", x"79787879",
									 -- x"7776787C", x"7D797879", x"7F7D7B7B", x"7C7C7F81", x"82828384", x"86868685", x"8A888888", x"87838180",
									 -- x"82828282", x"82827F7E", x"7C7D7C7A", x"7B7D7B77", x"78777776", x"75747678", x"7D7B7A7B", x"7E7F7F7D",
									 -- x"7D80817F", x"7E7F8182", x"83838283", x"85878888", x"8A8B8D8F", x"9194979A", x"9C9C9EA2", x"A5A8AAAC",
									 -- x"B1B2B4B8", x"BCBFC1C2", x"C4C7C9CA", x"C9C9CBCD", x"CACACBCB", x"CBCBCCCC", x"C9C9C6C3", x"C2C3C2BF",
									 -- x"C2C0C0C1", x"C3C2C2C3", x"C6C6C6C5", x"C4C5C6C7", x"CCCBCAC9", x"C9C9CACA", x"CACACAC9", x"C9C8C7C7",
									 -- x"C9CACACA", x"CCD0D1D0", x"D0CECBC7", x"C4C2C1C0", x"BEBFC2C3", x"C5C6C5C4", x"C4C7C6C8", x"C8C4C7C4",
									 -- x"C3C4C5C8", x"CBCCCBCA", x"CAC7C3BF", x"BCB8B4B2", x"B1AFACA9", x"A8A6A3A1", x"9E9D9B98", x"94918F8D",
									 -- x"8B8A8784", x"82827F7B", x"7875716F", x"6E6C6A6A", x"65626060", x"605E5D5D", x"5B595755", x"54535251",
									 -- x"53515152", x"53535353", x"54525153", x"55565758", x"56585959", x"57555351", x"5352514F", x"4F4F4D4A",
									 -- x"4A494949", x"47454547", x"44444341", x"3F3D3C3C", x"3D3C3A39", x"37363434", x"37373839", x"3837393D",
									 -- x"403F3F42", x"464A4C4C", x"51535351", x"4F4E4943", x"3D3D3A36", x"383D3C37", x"37393B3D", x"3D3E3E3E",
									 -- x"3F3A3532", x"33322E2A", x"2C2C2B29", x"27252626", x"26252422", x"22212121", x"2124231F", x"1B1C1F20",
									 -- x"201F1E1E", x"1E1E1D1C", x"1C19191B", x"1C1A1B1E", x"1A1A1B1C", x"1E1E1C1A", x"1C1B1B1D", x"1E1D1B19",
									 -- x"1B1B1B1A", x"1A191715", x"15191B1A", x"1B1D1A15", x"18181919", x"18161719", x"18181818", x"1A1C1C1A",
									 -- x"1C1A191A", x"1B1B1B19", x"1B1A1818", x"191A1B1A", x"1C1B1A1A", x"1A1A1A1A", x"1B1B1B1B", x"1C1C1C1B",
									 -- x"1A1A1A1A", x"1A191919", x"1D1C1A19", x"1A1B1B19", x"1A171618", x"1B1B1A1A", x"191A1B1C", x"1C1B1B1A",
									 -- x"1B1B1B1B", x"1D1E1C18", x"181B1C1A", x"191A1B1B", x"1A1A1A1A", x"1A1B1B1A", x"1C1E1F1D", x"1C1C1C1C",
									 -- x"1F1D1C1D", x"1E1F1E1D", x"201F1F1F", x"1F202020", x"1F202325", x"25232120", x"22222222", x"22222323",
									 -- x"24262727", x"2727292A", x"2C2B2928", x"28292A2A", x"2A2A2C2E", x"2D2A2C31", x"2F302E30", x"33323034",
									 -- x"716F726F", x"6E706D70", x"70716F6A", x"696D706F", x"726F6E71", x"73727272", x"74767778", x"78797A7A",
									 -- x"7473767B", x"7C79797B", x"7C7A797B", x"7D7E8285", x"8686888A", x"8C8D8D8C", x"8D8E8F8F", x"8C898A8D",
									 -- x"89898A8B", x"8C8B8885", x"82858480", x"7E7F7F7C", x"7C807F7A", x"787C7E7D", x"807C7A7C", x"80828280",
									 -- x"7F828483", x"83858788", x"88868587", x"8C8E8D8B", x"8C8D8E90", x"91949798", x"9B9C9FA1", x"A4A8ABAC",
									 -- x"AFB0B1B4", x"B8BCBEBF", x"C2C4C6C6", x"C5C3C4C5", x"C7C6C5C5", x"C7C8C7C6", x"C4C4C2C0", x"BFBEBDBB",
									 -- x"BCBBBCBD", x"BCBBBDBF", x"C3C3C2C1", x"C0BFC0C1", x"C2C3C3C3", x"C2C2C1C1", x"C4C4C4C4", x"C4C3C2C2",
									 -- x"C4C5C5C5", x"C7C9CACA", x"CBC9C7C4", x"C1BEBDBC", x"BCBDBFC2", x"C2C2C1C1", x"C2C4C0C3", x"C4C2C5C2",
									 -- x"C2C2C2C4", x"C6C7C6C5", x"C1C1BFBD", x"B9B6B3B1", x"AFACA9A6", x"A4A3A09F", x"9B9A9996", x"938E8B8A",
									 -- x"8786837F", x"7D7B7774", x"72706D6A", x"69686664", x"625F5C5C", x"5B5A5858", x"58565452", x"504F4E4D",
									 -- x"504F4F52", x"54535455", x"58545255", x"595A5858", x"56585B5C", x"5B595756", x"54575957", x"55545251",
									 -- x"514F4D4E", x"4E4C4B4B", x"4B4D4C48", x"44424446", x"40414140", x"3F3D3C3B", x"3D404444", x"403B3C3F",
									 -- x"42424448", x"4C4F5051", x"585C5D58", x"54514D49", x"43423E3C", x"3F444542", x"40414445", x"45454545",
									 -- x"45454441", x"3B363332", x"33302D2A", x"29292828", x"27272523", x"22222323", x"25222021", x"201F2023",
									 -- x"2422201F", x"1F1E1D1D", x"1D1A191C", x"1C1A1A1D", x"1B1A1A1A", x"1C1C1B1A", x"1919191A", x"1B1C1B19",
									 -- x"1C1B1B1B", x"1B191716", x"17181713", x"14181A18", x"17161719", x"1816171A", x"16161617", x"191C1C1A",
									 -- x"18171719", x"1A1B1918", x"1B191818", x"191A1A1A", x"1C1A1918", x"191A1919", x"18191A1B", x"1B1A1919",
									 -- x"1A1A1919", x"1A1A1919", x"1A1A1A1A", x"1A191919", x"1B181618", x"1B1A1A1A", x"19191A1B", x"1B1A1A19",
									 -- x"1A1A1A1A", x"1C1D1B17", x"181A1C1B", x"1A1A1A1A", x"1A191818", x"18191A1B", x"1A1D1E1C", x"1B1B1C1C",
									 -- x"1C1B1B1C", x"1D1F1F1E", x"1F1E1D1C", x"1C1C1D1D", x"1E202224", x"25242220", x"1F202020", x"20202123",
									 -- x"23242525", x"25262729", x"2A292928", x"27282A2C", x"2B29292C", x"2C2B2C30", x"31312E2F", x"34333235",
									 -- x"73717470", x"6F706D70", x"6F70706F", x"6D6E6F6F", x"736E6B6E", x"71717171", x"6F727576", x"76777777",
									 -- x"75757779", x"78767677", x"7978797B", x"7B7C7F82", x"87888A8C", x"8E909191", x"95989A98", x"95969CA1",
									 -- x"99989899", x"9995908C", x"8A8B8984", x"807F7F7E", x"8084827C", x"7B80827F", x"817D7B7D", x"81838483",
									 -- x"83868786", x"86888A8A", x"8C8B8B8F", x"94979693", x"96969696", x"97999A9B", x"999B9D9F", x"A1A6A9AA",
									 -- x"ADAFB0B1", x"B5B9BBBB", x"BBBDC0C1", x"C1C1C1C2", x"C3C2C0C1", x"C3C4C2C0", x"BEBDBCBA", x"BAB9B7B6",
									 -- x"B7B7B9B9", x"B8B7B9BC", x"BCBDBEBE", x"BDBBBAB9", x"BBBBBCBD", x"BDBCBBBA", x"BCBCBDBE", x"BEBEBEBE",
									 -- x"BFBFBFC0", x"C0C2C2C3", x"C6C4C3C2", x"C0BDBBBC", x"BDBCBDBD", x"BDBBBCBE", x"BFC0BBBE", x"BFBEC2BF",
									 -- x"C1C0C0C0", x"C1C2C1BF", x"BCBDBDB9", x"B5B2AFAC", x"ABA9A7A4", x"A19F9E9C", x"97959493", x"918D8987",
									 -- x"82827F7B", x"7876726F", x"6E6C6864", x"6362605C", x"5E5A5857", x"57545353", x"5453514F", x"4E4D4C4C",
									 -- x"4E4B4B4E", x"51515356", x"5C585659", x"5D5E5C5B", x"5C5D5F61", x"615F5D5D", x"5A5E6160", x"5C5B5A59",
									 -- x"58555455", x"56545252", x"5154544F", x"4A494B4E", x"484A4A47", x"45454442", x"45494C4C", x"46414043",
									 -- x"41454B4E", x"4F4F5459", x"5B61625B", x"5553504B", x"45434244", x"484C4E4E", x"4A4C4E4F", x"50504F4E",
									 -- x"504E4E4F", x"4D463F3A", x"37353230", x"2F2D2927", x"27272624", x"22222324", x"29232023", x"25232326",
									 -- x"28252321", x"1F1D1C1D", x"1F1E1D1D", x"1C1B1A1B", x"1B1A1919", x"1A1A1A1A", x"18191919", x"1A1C1B1A",
									 -- x"1A19191A", x"1B1A1919", x"18171614", x"1417191A", x"16161718", x"17161719", x"15161717", x"191B1C1A",
									 -- x"1718181A", x"1B1A1918", x"19181819", x"1A1B1A19", x"19181818", x"191A1A1A", x"1A1B1C1D", x"1C1B1A1A",
									 -- x"1A191919", x"1A1A1919", x"1717191A", x"1918191A", x"1B19181A", x"1B1A1919", x"19191A1A", x"1A191918",
									 -- x"1A1B1B19", x"191B1915", x"1718191A", x"19191818", x"1B191717", x"1718191C", x"191A1B1A", x"1A1B1C1C",
									 -- x"19191A1A", x"1B1C1D1E", x"1F1F1D1C", x"1C1C1D1D", x"2020201F", x"21232322", x"20202121", x"20212223",
									 -- x"23242424", x"24242628", x"27282827", x"27282A2C", x"2B29282A", x"2B2B2C2E", x"2F2F2C2D", x"302F2F33",
									 -- x"78767975", x"74747173", x"71707071", x"706F6E6E", x"706B6A6E", x"716F6E6F", x"6E737777", x"76777775",
									 -- x"75777877", x"75757574", x"797A7D7E", x"7D7C7E81", x"8587898B", x"8E909294", x"9CA2A4A1", x"9FA3A8AA",
									 -- x"A6A6A6A6", x"A6A29B96", x"95928E8B", x"88858485", x"86868481", x"80838482", x"87828082", x"85868585",
									 -- x"888A8A89", x"8A8C8D8D", x"90929598", x"9C9D9D9D", x"A1A09F9F", x"A0A2A3A3", x"9C9FA09F", x"A0A4A6A7",
									 -- x"ABADAFB0", x"B3B6B7B5", x"B5B7B9BC", x"BEBEBEBD", x"BCBBBBBC", x"BDBCBBB9", x"B7B7B6B5", x"B5B4B2B1",
									 -- x"B4B3B4B5", x"B5B4B5B7", x"B5B6B8B8", x"B6B5B4B3", x"B4B5B6B7", x"B7B6B5B5", x"B3B4B4B5", x"B6B7B7B8",
									 -- x"B7B7B8B9", x"B9B9BABB", x"BEBCBCBD", x"BDBAB9BA", x"B9B8B9B9", x"B8B6B6B8", x"B9BBB8BA", x"BAB8BDBC",
									 -- x"BEBDBCBC", x"BDBCBBB9", x"B9BAB9B3", x"AEACAAA8", x"A6A5A3A1", x"9D9A9998", x"938F8D8D", x"8C888483",
									 -- x"7B7B7A76", x"74726F6C", x"6B68635F", x"5E5F5D59", x"5A565454", x"53514F4F", x"4F4E4C4B", x"4A4A4949",
									 -- x"4B494A4F", x"52525457", x"5C5B5C60", x"63656667", x"6867676A", x"6B6A6867", x"65686968", x"66656463",
									 -- x"605E5D5D", x"5C5A5858", x"585A5956", x"54545454", x"5354524D", x"4A4A4A49", x"4E4E4D4B", x"48444547",
									 -- x"474A4F53", x"5353575D", x"5E63635D", x"59595651", x"4A484B51", x"5657595C", x"5757595B", x"5D5D5B5A",
									 -- x"5D565255", x"58554D46", x"3D3C3A37", x"332F2B29", x"29282725", x"23222324", x"28252323", x"25262626",
									 -- x"27252423", x"211E1D1F", x"1F1F1F1D", x"1C1C1B19", x"1A1A1A19", x"18181919", x"18191A1A", x"1A1C1B19",
									 -- x"18161618", x"19181819", x"1616181A", x"19171616", x"16171716", x"14151718", x"14161717", x"17191A19",
									 -- x"19191A1A", x"1A191919", x"17171819", x"1B1B1917", x"18181919", x"19191919", x"1C1D1D1C", x"1B1A1B1B",
									 -- x"1A191819", x"1A1A1918", x"18171719", x"1918191A", x"1B1A1A1B", x"1B191819", x"1A1A1A19", x"19191818",
									 -- x"181B1B18", x"17191815", x"16161617", x"17171615", x"1A181617", x"1717181B", x"18181817", x"191B1C1A",
									 -- x"191A1A1A", x"18191B1D", x"1E1D1D1D", x"1D1D1D1D", x"1F1F1D1C", x"1D20211F", x"21202020", x"20202020",
									 -- x"23232423", x"22232527", x"28272626", x"27282828", x"292A2B29", x"282A2B2B", x"292A2929", x"2C2B2A2E",
									 -- x"7E7C7F7B", x"797A7678", x"77716E6F", x"706D6C6D", x"6A67696E", x"706E6C6E", x"696E7272", x"7171706E",
									 -- x"70747674", x"75787A79", x"7A7D8184", x"84838588", x"8587898C", x"8E919496", x"9DA4A8A5", x"A4A8A9A6",
									 -- x"A7A7A9AB", x"ADABA5A0", x"A0999494", x"93908F90", x"8E8A8787", x"88878688", x"8D898788", x"89888686",
									 -- x"8A8B8C8C", x"8F939595", x"92969C9F", x"A0A1A2A4", x"A5A5A4A5", x"A6A8A9A9", x"A5A7A7A4", x"A3A5A7A7",
									 -- x"A9ACAEAF", x"B1B4B3B1", x"B6B6B8B9", x"BAB9B6B5", x"B4B6B7B7", x"B6B5B4B4", x"B4B3B3B3", x"B3B1B0AF",
									 -- x"B1AEADAF", x"B1B1B1B1", x"B2B2B1B0", x"AFAEAFB0", x"AEAFB0B1", x"B1B1B0B0", x"AEAEAEAF", x"AFB0B0B1",
									 -- x"B1B1B2B3", x"B3B3B4B6", x"B4B2B3B6", x"B6B4B3B4", x"B2B2B5B8", x"B6B3B1B2", x"B3B8B6B8", x"B6B3B9B9",
									 -- x"B8B8B7B7", x"B8B7B4B2", x"B1B3B1AC", x"A8A8A8A7", x"A1A1A09D", x"99959493", x"8F8A8685", x"85817D7C",
									 -- x"73747371", x"6F6E6C69", x"6966605C", x"5C5E5D5A", x"57545252", x"52504E4D", x"4B4A4847", x"46464545",
									 -- x"4A494E56", x"5A59585A", x"5B5D6166", x"696C7073", x"74707072", x"74737170", x"6F70706E", x"6E6E6D6B",
									 -- x"66656564", x"605C5B5C", x"5D5E5E5C", x"5C5E5C59", x"58585550", x"4D4E5051", x"534F4A47", x"4645474A",
									 -- x"52515256", x"595A5C5E", x"61656661", x"6062605A", x"514F545E", x"62606267", x"60606164", x"67676562",
									 -- x"625D5958", x"57555455", x"4443403B", x"35302E2D", x"2A2A2926", x"24222324", x"25262522", x"23272724",
									 -- x"25242424", x"23201F21", x"1C1F1E1B", x"1B1C1B18", x"191A1A19", x"17171719", x"16181919", x"191A1816",
									 -- x"18161517", x"17161617", x"17151619", x"18141315", x"16181814", x"13151716", x"13161716", x"15161717",
									 -- x"18191918", x"16151618", x"1616171A", x"1B1A1816", x"18191A1A", x"19181818", x"1B1B1A18", x"17161819",
									 -- x"1A191818", x"1A1A1918", x"1C181617", x"19191819", x"1B1A1B1C", x"1B191819", x"1B1B1A19", x"19181818",
									 -- x"161A1A17", x"16191917", x"19171616", x"17181717", x"19171618", x"18171719", x"17171615", x"171A1B19",
									 -- x"1A1C1C1A", x"18171A1C", x"191A1B1C", x"1C1C1B1B", x"1C1D1D1B", x"1D1F1E1B", x"1E1D1C1B", x"1C1C1B1A",
									 -- x"23232323", x"22222426", x"29272425", x"27282624", x"252B2D29", x"27282A29", x"25282829", x"2C2A2A2E",
									 -- x"8A8B8A87", x"8688847E", x"7F797270", x"7273716E", x"6B686769", x"6B6B6B6C", x"676B6E6E", x"6F6F6D69",
									 -- x"72737373", x"73757A7E", x"80848788", x"888A8B8B", x"8D898788", x"8C909599", x"9D9EA2A8", x"A8A5A6A9",
									 -- x"A6A7A9AB", x"ADACA8A5", x"A5A29F9C", x"9B999795", x"92908F90", x"91918D8A", x"8E909292", x"908E8D8D",
									 -- x"8A8D9093", x"96999C9E", x"9E9DA0A6", x"A7A5A6A9", x"ABABADB1", x"B2B1B1B2", x"B2B0ADAA", x"A8A6A5A5",
									 -- x"A9ABAEB0", x"B3B5B4B1", x"B4B6B7B5", x"B4B5B5B4", x"B1B3B3B1", x"B0B1B0AE", x"ADAEAEAD", x"ABAAAAAB",
									 -- x"ACAAA9A8", x"A8A8A8A8", x"A9A9A9A9", x"A9A8A7A7", x"A9A9AAA9", x"A8A7A8AA", x"A7A8A8A9", x"A9A9A8A8",
									 -- x"A9ABABAA", x"ABACABA9", x"AEAEAEAF", x"B0B0B0B0", x"B1B2B4B4", x"B2B1B1B1", x"B4B2B1B1", x"B1B2B2B2",
									 -- x"B4B0AEB0", x"B1AFACAA", x"A8A8A8A7", x"A5A3A09F", x"9F9D9A97", x"93908D8B", x"89868380", x"7D7B7875",
									 -- x"736F6D6D", x"6D696563", x"655F5B5C", x"5C5A5858", x"53535151", x"504E4C4B", x"4946474A", x"4A464445",
									 -- x"494C4E53", x"595A595D", x"61656768", x"6C74797B", x"81828683", x"7E7D7A7D", x"7679797A", x"77767B76",
									 -- x"716F6D6B", x"68646262", x"62606060", x"6064645F", x"53595B57", x"53545453", x"5A544E4C", x"4D4E4F51",
									 -- x"5757585A", x"5D606466", x"6864656D", x"6F69615E", x"5B5B5C5F", x"64696C6E", x"6C6D6E6F", x"6F6F6D6B",
									 -- x"67676663", x"605D5B5A", x"514A423E", x"3B363130", x"2B2C2A27", x"25252320", x"22212123", x"25252321",
									 -- x"22201F21", x"22222122", x"1C1C1C1C", x"1B1B1A1A", x"161B1C18", x"15171716", x"18151519", x"1814151A",
									 -- x"1C181516", x"16141314", x"13151617", x"16161515", x"16141213", x"15151412", x"16161515", x"15151616",
									 -- x"14171716", x"15161615", x"15161616", x"17171819", x"18191A1B", x"1B1A1817", x"191A1B1A", x"1818191A",
									 -- x"1D1C1A19", x"19191817", x"1517191A", x"19181717", x"1A191818", x"19191918", x"18181818", x"18181818",
									 -- x"15141415", x"16171514", x"16161616", x"15151414", x"17161515", x"16161616", x"17151415", x"17181817",
									 -- x"1C1B1917", x"16161718", x"1B1D1D1C", x"1A181819", x"1A1B1B1A", x"1A1D1E1E", x"1D1C1D1E", x"1D1C1D1F",
									 -- x"1F212426", x"25232427", x"25252627", x"26242426", x"2A272527", x"29272627", x"27292A2A", x"2D2F2F2E",
									 -- x"999B9A97", x"9696918A", x"87837D79", x"7775716F", x"6C69696A", x"6B6A6969", x"67696A6A", x"6B6D6D6B",
									 -- x"6E707171", x"7073797E", x"81838483", x"83858889", x"8C898887", x"888A8F94", x"9B9A9EA4", x"A5A3A3A5",
									 -- x"A1A1A2A5", x"A9ACACAB", x"A7A5A3A2", x"A3A2A09E", x"9B999796", x"9493908E", x"92949696", x"94939293",
									 -- x"91939697", x"9A9DA2A6", x"ABA9A7A8", x"A9ABAFB3", x"B5B4B3B2", x"B3B4B4B4", x"B0AFACAA", x"A7A7A7A8",
									 -- x"A8AAACAE", x"B0B3B2B0", x"B2B3B2AF", x"AEAFAFAE", x"AAABAAA8", x"A8AAAAA8", x"A7A7A8A7", x"A5A4A3A4",
									 -- x"A2A1A0A0", x"A0A1A1A0", x"A1A1A1A0", x"A09F9F9E", x"A1A1A2A1", x"A09FA0A0", x"9F9E9E9F", x"9FA0A1A1",
									 -- x"A3A4A4A3", x"A4A6A5A2", x"A6A6A6A7", x"A8A8A8A8", x"A8AAABAC", x"ABABABAC", x"ADABAAA9", x"AAABACAC",
									 -- x"ACAAAAAB", x"ABA9A8A8", x"A6A6A5A3", x"A09D9A98", x"99979592", x"908D8B89", x"84827F7C", x"7A787573",
									 -- x"726F6B6A", x"68656160", x"605B5656", x"56555454", x"51504E4D", x"4C4C4B4B", x"4946474A", x"4A474547",
									 -- x"464A4D53", x"5B5C5D61", x"636A7174", x"767B8388", x"97959190", x"908E8C8A", x"8A857F85", x"8A898678",
									 -- x"7A75716E", x"6C686767", x"65636363", x"62656762", x"5C60615C", x"59595855", x"5D545258", x"58525259",
									 -- x"5B5C5E60", x"63676A6D", x"746F6C6F", x"716E6A69", x"66646363", x"666B7074", x"75757677", x"77757270",
									 -- x"68696967", x"65646465", x"61584E47", x"413A3431", x"2D2D2B27", x"25252422", x"22212223", x"25252322",
									 -- x"211F1E20", x"21212021", x"1C1C1B1A", x"19181818", x"14181915", x"13151614", x"18161618", x"17141518",
									 -- x"16131213", x"15151619", x"13141515", x"15151516", x"15151414", x"14141313", x"12131415", x"15151414",
									 -- x"14161715", x"15161615", x"15161615", x"15151616", x"18171615", x"15161718", x"17191A19", x"1817191A",
									 -- x"19181717", x"18181716", x"17171716", x"16161717", x"17171818", x"18181717", x"18181817", x"16151313",
									 -- x"15151312", x"12131517", x"16161615", x"15151515", x"16151414", x"14151616", x"15141414", x"16161514",
									 -- x"19181716", x"16161617", x"1A1A191A", x"1A1A1A1A", x"1B1D1E1E", x"1D1E1C1A", x"1C1C1C1D", x"1C1B1C1E",
									 -- x"22222325", x"24222224", x"27262526", x"25242526", x"2727292C", x"2B292828", x"292B2C2A", x"2A2C2D2E",
									 -- x"A5A7A7A4", x"A2A19B95", x"8E8B8782", x"7F7C7978", x"73716F6E", x"6C6A6969", x"67676766", x"686A6C6C",
									 -- x"696C6E6E", x"6D70767C", x"7B7D7D7D", x"7E83898C", x"8B898887", x"86868A8F", x"9291949B", x"9E9E9FA1",
									 -- x"9E9E9FA1", x"A5A8A9A9", x"A9A8A8AA", x"ADAEACAA", x"A5A4A29F", x"9C9A9898", x"9A9B9C9C", x"9C9A9A9A",
									 -- x"999C9EA0", x"A2A6ADB2", x"B4B2AEAA", x"AAAEB3B5", x"B9BAB8B5", x"B5B7B5B2", x"ADACABA8", x"A7A7A8A9",
									 -- x"A5A6A7A9", x"ACB0B0AF", x"AEADAAA7", x"A5A6A7A6", x"A5A5A4A2", x"A2A3A4A3", x"A0A1A1A1", x"9F9E9D9D",
									 -- x"9A999999", x"99999998", x"99999998", x"97979696", x"97989898", x"98989898", x"98979796", x"97979899",
									 -- x"9A9B9A9A", x"9B9C9B9A", x"9D9E9E9F", x"9FA0A0A0", x"9FA1A3A4", x"A4A5A5A6", x"A5A4A3A2", x"A3A4A5A6",
									 -- x"A3A3A4A4", x"A3A0A1A2", x"9F9F9F9E", x"9C999795", x"92908E8C", x"8B898785", x"827F7B78", x"75726F6D",
									 -- x"706B6866", x"64605E5D", x"5C585453", x"53525151", x"504F4C4B", x"4B4B4B4B", x"49464649", x"4A474748",
									 -- x"494C4F54", x"5B5C5C60", x"676D777E", x"81868D94", x"999D9AA6", x"AEACACA2", x"9E9C999D", x"9C97958C",
									 -- x"867F7773", x"706E6C6C", x"68666665", x"62646663", x"61646360", x"5D5D5A56", x"5854565C", x"5B555459",
									 -- x"57595D62", x"676C7072", x"7A777474", x"76777675", x"72706C69", x"696E757A", x"7D7B7875", x"736F6C6B",
									 -- x"6C6D6C69", x"66656668", x"6A61554C", x"443D3632", x"302F2C28", x"26262524", x"1E1E1E1F", x"1F1E1D1D",
									 -- x"1F1D1D1E", x"1F1F1F20", x"1C1B1A19", x"18171616", x"14181815", x"14151716", x"16171716", x"15141515",
									 -- x"17151413", x"13131619", x"14141313", x"13141617", x"15151615", x"13121314", x"11131517", x"17161413",
									 -- x"13151615", x"14151615", x"16171717", x"16161617", x"18171514", x"15161819", x"16171818", x"17171819",
									 -- x"16151515", x"16161515", x"16161514", x"14141515", x"13161819", x"18161515", x"18181918", x"17151311",
									 -- x"13141412", x"10111416", x"15151515", x"15151515", x"15141212", x"13141515", x"14141515", x"15141413",
									 -- x"16161717", x"17171717", x"19171617", x"1A1B1B1A", x"1C1E1F1E", x"1D1D1C1A", x"1C1B1C1D", x"1D1C1D1F",
									 -- x"221F1F20", x"21201F1F", x"26232222", x"22222325", x"2526292B", x"29272728", x"2A2D2E2C", x"2A2B2E2F",
									 -- x"A9AAA9A7", x"A6A5A29F", x"97928C87", x"83817E7D", x"7D7A7774", x"716E6D6C", x"67666565", x"66686868",
									 -- x"67686A6B", x"6B6E7275", x"74767777", x"7A808588", x"85838282", x"8284878B", x"8A898B90", x"94959595",
									 -- x"97989B9E", x"A2A4A5A5", x"A8A7A9AD", x"B1B3B1AF", x"AEADABA9", x"A7A5A4A3", x"A2A2A3A3", x"A3A19F9D",
									 -- x"9EA2A6A9", x"ABAEB4B9", x"B7B7B3AE", x"ADB1B2B0", x"B4BABBB7", x"B5B6B3AD", x"ACAAA8A7", x"A7A7A6A5",
									 -- x"A6A5A5A5", x"A8AAAAA9", x"A8A7A4A1", x"A0A0A1A0", x"A2A1A09F", x"9E9D9D9C", x"999A9B9B", x"9A989796",
									 -- x"96959494", x"93929190", x"93929291", x"9090908F", x"8D8E8E8F", x"8F909292", x"92929191", x"90909090",
									 -- x"92929292", x"93939392", x"95969797", x"98989898", x"98999A9C", x"9D9E9E9F", x"9E9D9D9D", x"9E9F9F9E",
									 -- x"9E9E9E9D", x"9B9A9A9A", x"97979796", x"95939190", x"8C8B8987", x"85838180", x"7D7A7673", x"716E6B69",
									 -- x"6A666362", x"605D5B5B", x"5B585554", x"53525150", x"51504E4D", x"4C4C4C4C", x"4C49494B", x"4C4A4A4C",
									 -- x"4C505256", x"5C5D5E63", x"6D727C86", x"8D92989D", x"A4AEABBA", x"C1BABEB3", x"AFB3B6BA", x"B2A6A298",
									 -- x"8D847A75", x"72706D6B", x"68666765", x"6160625F", x"5F605F5D", x"5C5C5955", x"50555854", x"53555653",
									 -- x"595B5F66", x"6E747676", x"76777879", x"7C7F7E7B", x"79787571", x"6F71767B", x"837E7771", x"6D6B6B6B",
									 -- x"6A6A6965", x"62606265", x"675F544B", x"443E3835", x"312F2B28", x"27262422", x"21222221", x"1F1E1D1E",
									 -- x"1D1B1B1C", x"1D1C1C1E", x"1C1B1918", x"17161616", x"14161614", x"13151616", x"14161613", x"13151513",
									 -- x"16161513", x"12111315", x"14141413", x"13131516", x"15151514", x"13131313", x"11131517", x"17161412",
									 -- x"13141414", x"14141516", x"15161617", x"16161717", x"16161718", x"18171717", x"15161716", x"16151617",
									 -- x"16151414", x"14141414", x"14141515", x"15141211", x"12151718", x"16141415", x"14151718", x"17161413",
									 -- x"11121313", x"12121213", x"14141414", x"13131313", x"13131212", x"13141515", x"15161616", x"15151516",
									 -- x"16161717", x"18181818", x"19181717", x"18191A1A", x"1B1C1C1A", x"1A1C1D1C", x"1C1C1C1E", x"1E1E1F21",
									 -- x"1F1D1C1E", x"1F1F1F20", x"24212021", x"22232324", x"25252525", x"24242527", x"272A2B2A", x"2A2C2E2F",
									 -- x"A9A9A7A6", x"A7A8A9A9", x"A79F948C", x"87847F7B", x"7E7F7F7D", x"7976726F", x"6B696868", x"68676564",
									 -- x"67666668", x"6B6D6D6C", x"6E717373", x"74787B7C", x"7B787679", x"7C7F8082", x"87868688", x"8A8A8988",
									 -- x"8A8C9095", x"9A9FA2A3", x"A4A5A8AD", x"B1B3B2B0", x"B4B1AFAE", x"AFAFADAB", x"A6A7A8AA", x"AAA8A5A2",
									 -- x"A3A8AEB1", x"B3B4B7B9", x"BABBB9B4", x"B3B5B3B0", x"B1B8BAB5", x"B1B0AFAB", x"ACA9A6A7", x"AAAAA6A2",
									 -- x"AAA8A6A5", x"A5A4A2A1", x"A3A19F9F", x"9F9E9D9C", x"9C9B9B9A", x"98959392", x"92929393", x"9391908E",
									 -- x"8F8E8D8D", x"8C8B8988", x"8B8A8988", x"88878787", x"86858484", x"8687898A", x"89898A8A", x"89898787",
									 -- x"8B8A8A8B", x"8B8B8B8B", x"8C8D8E8F", x"8F8F8F90", x"90919192", x"94949595", x"95959596", x"97979695",
									 -- x"97979695", x"95959493", x"9191908E", x"8C898786", x"88868482", x"7F7D7B79", x"7573716F", x"6E6C6A69",
									 -- x"6461605F", x"5E5A5959", x"5A595655", x"54535150", x"51505050", x"504F4F4E", x"504F4E4F", x"504F4F50",
									 -- x"4F525459", x"5F62656B", x"707B8B96", x"9B9EA5AB", x"B4C0BEC9", x"CBC7D3D0", x"CECBC8CF", x"CDC0AE96",
									 -- x"8C837975", x"73706C69", x"68666766", x"615E5E5B", x"5C5B5A58", x"58575451", x"4E53534E", x"4D515453",
									 -- x"5C5D6068", x"70747370", x"76797B7D", x"80817F7B", x"7B7C7B79", x"76747577", x"7C76706C", x"6967686A",
									 -- x"63636260", x"5D5D5F62", x"625D544C", x"45403C39", x"312E2B29", x"28252220", x"21212120", x"1E1D1D1D",
									 -- x"1C1A1A1B", x"1B191A1B", x"1A191816", x"15151516", x"11121312", x"11121313", x"12151512", x"12151512",
									 -- x"10121312", x"11121415", x"14141414", x"13131314", x"16141313", x"14141311", x"11121314", x"13121110",
									 -- x"12121313", x"13131415", x"13141515", x"14141415", x"13141516", x"16151312", x"15151515", x"14131414",
									 -- x"16151413", x"12131415", x"14141414", x"14141211", x"12141616", x"14131416", x"10111314", x"15141312",
									 -- x"12121112", x"13131211", x"12121212", x"12121212", x"13121314", x"15151414", x"16161615", x"15151617",
									 -- x"17161616", x"16171819", x"18181818", x"1717191A", x"1A1B1B1A", x"1A1C1D1C", x"1B1B1C1E", x"1E1E1F22",
									 -- x"1F1E1E20", x"201F2124", x"23222224", x"26252527", x"24242222", x"24252625", x"24262728", x"2A2C2C2A",
									 -- x"A4A3A3A2", x"A4A7AAAB", x"B0A89D96", x"928D8781", x"7D818586", x"837E7873", x"73706E6E", x"6E6A6663",
									 -- x"68666466", x"6A6C6966", x"696C6F70", x"70727474", x"74706F72", x"77797979", x"7E7E7F81", x"82838484",
									 -- x"82838589", x"8E94999C", x"A2A5A9AD", x"B1B2B3B3", x"B5B1AEAE", x"B1B2B1AF", x"ADADAFB1", x"B3B3AFAC",
									 -- x"ADB1B6BA", x"BBBABAB9", x"BEBDBAB7", x"B7B7B6B4", x"B4B7B7B1", x"ADADADAC", x"AAA7A5A6", x"AAABA7A2",
									 -- x"A7A5A4A5", x"A5A3A2A1", x"9F9D9C9D", x"9D9B9998", x"96959595", x"93908D8C", x"8D8D8D8D", x"8D8C8B89",
									 -- x"89888786", x"86858483", x"83838280", x"807F7F7F", x"81807E7E", x"7F808181", x"7E7F8182", x"8281807F",
									 -- x"84828182", x"83838383", x"84868787", x"87868789", x"8B8A8A8B", x"8C8C8C8C", x"8D8E8E8F", x"908F8E8D",
									 -- x"8D8D8C8B", x"8C8D8D8B", x"89898887", x"85848281", x"817F7D7B", x"79777473", x"73706D6B", x"6A686563",
									 -- x"615F5E5E", x"5C595758", x"59595856", x"55555452", x"53535354", x"55555453", x"54535253", x"54545454",
									 -- x"5558595C", x"6164676E", x"72879EA6", x"A5A7B2BC", x"BDC8CDD9", x"DDDFEBEC", x"EFE7D9D7", x"D6CEBC9F",
									 -- x"8C847C78", x"76726E6B", x"69656565", x"605C5B58", x"5B595654", x"53514F4D", x"4F4A4A4D", x"4D4A4F57",
									 -- x"5A5D636B", x"72757370", x"797A7C7D", x"7D7C7B7A", x"797B7B7A", x"78757473", x"736F6B6A", x"67625F60",
									 -- x"61615F5D", x"5B5A5A5B", x"5D5C564D", x"46413D3B", x"34302D2C", x"2A272321", x"1E1E1C1B", x"1B1B1B1B",
									 -- x"1B1A1A1A", x"19171719", x"17161514", x"13131313", x"11111212", x"12121211", x"12131311", x"11141412",
									 -- x"10121313", x"13141514", x"13141414", x"13121111", x"15131112", x"14141311", x"13131312", x"12111111",
									 -- x"13121212", x"12111315", x"14141515", x"14131212", x"14131313", x"12121212", x"14141313", x"13121211",
									 -- x"14141312", x"12131516", x"16141111", x"12131313", x"13131413", x"12121415", x"11111213", x"13121211",
									 -- x"15120F0F", x"10121212", x"11111111", x"11111112", x"13131314", x"15151413", x"15151414", x"15151516",
									 -- x"16151515", x"15161717", x"17181919", x"18181A1C", x"1A1C1D1D", x"1C1D1B19", x"1A1A1B1C", x"1D1C1E20",
									 -- x"1E1E1E1F", x"1F1E1F22", x"20212325", x"25242426", x"23232425", x"282A2826", x"2628292A", x"2C2E2C2A",
									 -- x"98999A9B", x"9C9EA0A1", x"A6A39F9C", x"9B97918C", x"858A8D8D", x"8A86817D", x"7E797675", x"736F6A68",
									 -- x"6A676465", x"686A6865", x"65686969", x"696C6E6F", x"6D6B6A6E", x"71737374", x"7476787A", x"7B7E8081",
									 -- x"7D7E7F82", x"85898E90", x"9B9FA5A9", x"ACADB0B1", x"B0ADAAAA", x"ACAFB1B2", x"B3B2B2B4", x"B8B8B6B3",
									 -- x"B4B6B9BC", x"BDBDBBBA", x"BDB9B7B7", x"B8B8B7B7", x"B5B4B2B0", x"AFAEADAD", x"A8A6A4A4", x"A5A5A4A2",
									 -- x"9E9D9EA2", x"A5A4A2A2", x"9E9B999A", x"9A979594", x"908F8F90", x"8F8C8A8B", x"89888888", x"88888685",
									 -- x"84838280", x"80807F7E", x"7D7C7B7A", x"79797979", x"7B7A7979", x"797A7978", x"76777879", x"7A7A7979",
									 -- x"7B787879", x"7A79797B", x"7C7D7F7F", x"7E7E7F81", x"84838283", x"84858584", x"87868686", x"86868584",
									 -- x"81838381", x"80828382", x"8080807F", x"7E7D7C7C", x"78777573", x"72706F6D", x"706D6A67", x"6663615E",
									 -- x"62605F5F", x"5D5B5C5D", x"5E5E5D5B", x"5B5D5D5C", x"5D5C5C5C", x"5D5D5D5C", x"5A5A5A5A", x"5B5C5C5C",
									 -- x"60626263", x"67696D75", x"8397A9AB", x"A9B0BFC9", x"D0D4D9E2", x"EAEDEDEB", x"F5F2E4DA", x"D2CCBDA3",
									 -- x"8E867E79", x"75716C6A", x"66605F5F", x"5B585855", x"5856524F", x"4D4B4949", x"4943454D", x"4F4B4E58",
									 -- x"5C636C73", x"75757575", x"76747678", x"78757578", x"76767574", x"73717070", x"716D6B6B", x"68625D5E",
									 -- x"605E5C5A", x"59575554", x"5758564E", x"45403E3C", x"3934302F", x"2D2A2625", x"2523201F", x"1F1F1E1D",
									 -- x"1B1A1A19", x"17151517", x"16161514", x"13121111", x"11111213", x"13121110", x"13121111", x"12121211",
									 -- x"14151412", x"12141412", x"11121312", x"11111010", x"13121112", x"13131211", x"14131312", x"12121213",
									 -- x"13121112", x"11101114", x"14151515", x"14131212", x"14131312", x"12121314", x"13121212", x"12111110",
									 -- x"12121312", x"12111213", x"15121010", x"11131312", x"12121111", x"11121313", x"14131212", x"11111111",
									 -- x"13110F0E", x"0E0F1111", x"10101111", x"12131313", x"15141312", x"13141414", x"15141415", x"16161412",
									 -- x"14141515", x"16161616", x"17181919", x"191A1B1B", x"1A1C1D1C", x"1C1C1A18", x"1C1B1B1C", x"1C1B1C1E",
									 -- x"1D1C1B1C", x"1D1D1D1E", x"1E1F2224", x"22202124", x"23252625", x"26282825", x"282A2C2C", x"2C2E2D2C",
									 -- x"8F909395", x"96969696", x"98999B9C", x"9B98928E", x"92949591", x"8D8B8986", x"86807A78", x"76726E6D",
									 -- x"6A676565", x"66676766", x"64656462", x"60626465", x"66656669", x"6C6D6F70", x"72747575", x"7677797B",
									 -- x"787A7D81", x"8486888A", x"90969DA1", x"A3A5A9AC", x"AAA8A6A5", x"A7ACB1B4", x"B4B2B0B2", x"B5B6B4B2",
									 -- x"B3B3B4B7", x"B9BAB9B8", x"BAB6B5B9", x"BBB9B8B9", x"B3B0AEB1", x"B3B1AEAC", x"A6A5A3A1", x"9F9E9F9F",
									 -- x"9C9A9CA0", x"A2A09E9E", x"9E9A9898", x"97949190", x"8B89898B", x"8B88888A", x"84838282", x"83828180",
									 -- x"82807E7C", x"7B7A7978", x"78777674", x"73737374", x"73737374", x"75747271", x"71717172", x"72727272",
									 -- x"74727173", x"73727374", x"73757777", x"76767779", x"7D7C7B7B", x"7D7E7D7D", x"807F7D7C", x"7D7D7D7D",
									 -- x"797D7D7A", x"77787A7B", x"7A7A7977", x"75747271", x"71706F6E", x"6D6C6B6A", x"68676564", x"64636261",
									 -- x"63616060", x"60606164", x"65666461", x"61656868", x"69676564", x"64646463", x"62626364", x"65676766",
									 -- x"696B6A6C", x"71747982", x"99A5ACA9", x"ABBAC9D0", x"DFD7D8DD", x"E9F2EDE9", x"E5E8E2DB", x"D3C9B492",
									 -- x"8D857C76", x"706B6664", x"625A5758", x"55545452", x"54514E4B", x"48464546", x"4243474D", x"51525457",
									 -- x"5A636D71", x"6D69696B", x"6D6B6E73", x"74707176", x"74726F6D", x"6D6D6D6D", x"66636163", x"625E5C5E",
									 -- x"5A585757", x"58575553", x"5156564F", x"46424040", x"3E383231", x"302C2928", x"2724201E", x"1E1D1B1A",
									 -- x"1B1A1A19", x"17141416", x"17171615", x"13121110", x"0F0F1011", x"12100E0D", x"14121011", x"12111010",
									 -- x"11110F0E", x"0F12120F", x"10111110", x"100F1010", x"11111212", x"11111213", x"11111110", x"11111112",
									 -- x"13111112", x"11101114", x"10121313", x"12111111", x"11111212", x"12121212", x"12111111", x"11111110",
									 -- x"11121313", x"110F0F0F", x"12111011", x"13131210", x"11101010", x"11121211", x"1312100F", x"0E0E0F10",
									 -- x"0E101111", x"0F0E0E0F", x"0F0F1011", x"13141515", x"16141211", x"11121414", x"15141517", x"18171310",
									 -- x"13141617", x"18181717", x"1A191819", x"1B1C1B19", x"1A1B1A18", x"181A1A19", x"1E1D1D1D", x"1C1A1B1D",
									 -- x"1E1B191C", x"1F1F1D1D", x"1F212324", x"211E2024", x"24262622", x"21222425", x"25292B2A", x"292B2C2D",
									 -- x"898B8E8E", x"8C8A898A", x"8E8D9096", x"98969494", x"9696938F", x"8E8F8F8D", x"868A887E", x"7977726B",
									 -- x"6D6C6B69", x"6A6B6964", x"6163625E", x"5C5D5F5F", x"61616367", x"696B6E72", x"6F727473", x"74757574",
									 -- x"73767A7C", x"7B7C848D", x"8A939B9F", x"A0A1A4A6", x"A3A5A3A0", x"A2A9ABAA", x"AAABAAAC", x"AEADADB2",
									 -- x"AFB1B3B4", x"B5B6B4B1", x"B5B3B2B5", x"B6B5B5B5", x"ADADAFB0", x"AEAAA9AB", x"A5A6A6A2", x"9D9A9B9E",
									 -- x"9A999898", x"9A9A9A99", x"96989995", x"908E8E90", x"8787888B", x"8A878483", x"84838383", x"8484817D",
									 -- x"7C7A7979", x"79787470", x"72717473", x"6E6C6D6B", x"696D6B6F", x"706E706C", x"6E6E6D6D", x"6E6F7071",
									 -- x"6F6F6D6B", x"6A6C6D6C", x"6C6E7070", x"70707173", x"75757576", x"77777878", x"78757476", x"76747373",
									 -- x"73737373", x"73737372", x"716F6E6F", x"6F6F6D6B", x"6E6C6A68", x"68686969", x"66636163", x"65625E5C",
									 -- x"61656869", x"68686A6C", x"706F6963", x"646C7375", x"75787471", x"76757173", x"76757573", x"72767771",
									 -- x"7675787B", x"7C859196", x"A6ADB5AE", x"AEC1CED4", x"E6DDD9E6", x"FAFCF2EB", x"EDEBDBCF", x"CCC4AC8A",
									 -- x"81797572", x"6A656361", x"5D595654", x"5154544F", x"4D4B4C4A", x"43404242", x"4040454C", x"5255575A",
									 -- x"60666E71", x"6C656262", x"62666B6E", x"6F6E6D6C", x"706E6A66", x"65676867", x"62616162", x"615C5958",
									 -- x"58565351", x"50515253", x"5254524E", x"49443E39", x"3B393532", x"2F2E2C2B", x"27242221", x"201E1C1C",
									 -- x"191A1A19", x"17141414", x"13131312", x"11111213", x"0F101011", x"1111100F", x"11121211", x"10101011",
									 -- x"10101010", x"11100F0E", x"100F0F11", x"110F0F11", x"14110F0F", x"11131312", x"100F0F0F", x"10111111",
									 -- x"12100E0E", x"0E101111", x"13110F0F", x"0F0F0F0E", x"10101112", x"11101011", x"10111213", x"1311100F",
									 -- x"0D0E1011", x"110F0E0D", x"0E10110F", x"10121311", x"10101010", x"10100F0F", x"10101010", x"1111100F",
									 -- x"1012110F", x"0F111211", x"12100F11", x"14161514", x"11111213", x"14141414", x"10111214", x"15151312",
									 -- x"14151617", x"17161413", x"1717181A", x"19161617", x"1B1A1818", x"1A1B1B1B", x"191A1B1B", x"1B1B1C1C",
									 -- x"191B1E21", x"21222121", x"23212021", x"201F2124", x"28252321", x"22232424", x"26262626", x"27292C2F",
									 -- x"89878382", x"8285898C", x"89898B8F", x"918F8E8F", x"9393918F", x"8E8E8D8B", x"8B8C8C87", x"807A7573",
									 -- x"736F6B68", x"6969655F", x"5C5E5E5B", x"595A5C5C", x"5D5D6064", x"66676A6D", x"6C6E706F", x"6F717271",
									 -- x"73747777", x"76767C83", x"888F9698", x"98999A9A", x"9B9D9D9A", x"9BA0A2A1", x"A2A4A3A5", x"A8A7A6AB",
									 -- x"ABABABAB", x"ACAEAFAE", x"B0AEAEB0", x"B1AFADAD", x"ABABABAA", x"A7A6A6A6", x"A3A2A19F", x"9D9B9B9B",
									 -- x"99989797", x"97979695", x"94949391", x"8E8D8D8D", x"8D8B8989", x"8783807F", x"85858584", x"83817F7E",
									 -- x"7A797775", x"74757575", x"78767572", x"6B6A6C6A", x"696D6C6E", x"6D6A6D6A", x"696A6B6C", x"6C6B6968",
									 -- x"6B6B6865", x"62626260", x"68696A6A", x"6969696A", x"6B6D6E6F", x"70707071", x"726E6C6F", x"71706F6E",
									 -- x"6D6C6A69", x"69696969", x"68676667", x"68696867", x"69696968", x"68686869", x"67646364", x"65646362",
									 -- x"66696B6C", x"6C6E7275", x"76726D6C", x"6D727A80", x"898A8682", x"85878788", x"8A8A8D8C", x"87868A8D",
									 -- x"8C88898E", x"939DA5A5", x"A8ACB4B1", x"B3BEC9D8", x"E2DFDFE9", x"F7FAF6F7", x"F5E9D5CD", x"C0AA9A8C",
									 -- x"7D746F6C", x"6663615E", x"5C595754", x"50504F49", x"4B464544", x"403F4242", x"3F42474C", x"50555C63",
									 -- x"64676C6C", x"67615F61", x"5E616568", x"68686766", x"6A696663", x"62646463", x"615E5B5B", x"5A575656",
									 -- x"54535150", x"50515150", x"4E4F4E4A", x"4744413D", x"3C3A3632", x"302D2B2A", x"26242221", x"201D1C1C",
									 -- x"18191817", x"15141415", x"15141312", x"12121212", x"0E0F1011", x"11100E0D", x"0F0F0F0F", x"10101111",
									 -- x"10101010", x"10100F0E", x"0F0E0E10", x"100F0F11", x"0F0F0F0F", x"0F0F1010", x"10101010", x"10100F0F",
									 -- x"11100F0F", x"10100F0F", x"11100F0E", x"0F0F0F0E", x"0E0E0F10", x"0F0F1010", x"0F0F0F0F", x"0F0E0D0D",
									 -- x"0F0F0E0E", x"0E0E0E0F", x"0D0F0F0E", x"0F111210", x"11111010", x"0F101010", x"11100F0F", x"10101010",
									 -- x"0E0F0F0D", x"0E101110", x"12121112", x"13131312", x"13131313", x"14151616", x"11111213", x"13131110",
									 -- x"10111416", x"17171716", x"15141517", x"16131214", x"1A191819", x"1A1B1B1B", x"1A1B1B1B", x"1A1A1A1A",
									 -- x"18191C1D", x"1D1D1D1D", x"1E1D1E20", x"201F2123", x"25242323", x"24252525", x"26282A2B", x"2B2A2A2B",
									 -- x"82807F7F", x"82848584", x"85858789", x"89898A8B", x"8F908F8E", x"8E8E8D8A", x"8C8C8D8C", x"847B787B",
									 -- x"78736C68", x"6868635D", x"57585755", x"53545657", x"55565A5F", x"62646769", x"696B6C6C", x"6D6F7070",
									 -- x"72737475", x"75767A7F", x"83888E90", x"92939393", x"93979896", x"95989A9A", x"9B9E9E9F", x"A2A09EA2",
									 -- x"A4A5A5A4", x"A5A8AAAA", x"A9A8A8AB", x"ABAAA7A6", x"A6A8A7A3", x"A2A4A6A4", x"9F9C9A99", x"99989693",
									 -- x"93929191", x"9292918F", x"91908E8C", x"8B8A8989", x"8A888788", x"86838182", x"83848584", x"817E7E7E",
									 -- x"7A787573", x"7173777A", x"79787876", x"6E6A6864", x"666B696B", x"69656968", x"65666768", x"67656361",
									 -- x"64646360", x"5F60605F", x"61626262", x"61616162", x"61646667", x"67666769", x"6A676466", x"69696766",
									 -- x"67656361", x"60606161", x"65656565", x"67696A6A", x"6D6E6F6F", x"6D6C6C6C", x"68666465", x"66656667",
									 -- x"6C6F7274", x"75777A7D", x"7D787576", x"7779818A", x"97969592", x"8E919493", x"95979995", x"92949A9F",
									 -- x"9D9A9DA4", x"ABB5BCBB", x"BAB6B6B9", x"C1C5CADD", x"E5E4E4EA", x"F4F9FBFF", x"FFEDD8CF", x"BC9E8E87",
									 -- x"7C726C69", x"6563625D", x"5B595854", x"4E4B4A44", x"48413F41", x"40424646", x"42474E52", x"53566069",
									 -- x"67686866", x"605B5B5E", x"5A5C5F61", x"61616161", x"61615F5D", x"5D5E5E5C", x"5B585554", x"53515151",
									 -- x"504F4E4E", x"4D4C4B4A", x"48494846", x"45444240", x"3E3C3834", x"312F2C2B", x"26232121", x"1F1D1B1B",
									 -- x"1A1A1817", x"15141415", x"16151312", x"12121110", x"0E0F1011", x"100F0D0B", x"110F0E0E", x"0E0E0D0C",
									 -- x"0F0F0F0F", x"0F0F0E0D", x"0D0D0D0E", x"0F0E0F10", x"0E0F1010", x"0F0E0E0F", x"0E101010", x"0E0E0E0F",
									 -- x"0F0F0F10", x"11100F0D", x"0F0E0D0D", x"0E0E0E0D", x"0C0C0D0D", x"0D0D0E0F", x"0F0F0E0E", x"0D0C0C0C",
									 -- x"0E0E0D0D", x"0D0D0E0E", x"0C0E0E0D", x"0E0F100F", x"100F0E0E", x"0E0F1011", x"11100F0E", x"0F101010",
									 -- x"0F10100F", x"0F111110", x"11121313", x"12111112", x"14131313", x"13141516", x"14131314", x"14131211",
									 -- x"12131414", x"15151414", x"18171818", x"17151517", x"17161617", x"18181818", x"18191919", x"18181819",
									 -- x"191A1C1C", x"1C1C1C1D", x"1C1C1E20", x"20202122", x"23232325", x"26272625", x"27292B2D", x"2C2B2A29",
									 -- x"7D7D7E80", x"81807D7A", x"7F808181", x"82828486", x"8A8A8A8A", x"8B8C8B8A", x"88878887", x"827C7A7B",
									 -- x"79746D6A", x"69686460", x"56555350", x"4F505254", x"5052565A", x"5D606264", x"64666869", x"6A6B6C6C",
									 -- x"6E6F7073", x"76797D7F", x"7F828587", x"8A8D8E8D", x"8C909291", x"90929494", x"95999999", x"9B999698",
									 -- x"9B9EA0A0", x"A1A2A2A1", x"A2A1A2A3", x"A5A5A4A3", x"A2A5A49E", x"9DA0A09D", x"9A979492", x"92908C89",
									 -- x"89888889", x"8B8B8A89", x"8E8D8C8C", x"8A888787", x"83838587", x"87848384", x"80818384", x"827F7E7F",
									 -- x"79787674", x"7475787A", x"7A777875", x"6E6A6864", x"64666467", x"66636767", x"66656362", x"61606061",
									 -- x"6060605E", x"5E616262", x"5C5C5C5C", x"5D5D5E5E", x"5B5E6060", x"5E5E6062", x"64615F5F", x"60605F5E",
									 -- x"6261605E", x"5D5D5E5F", x"63646566", x"686B6D6F", x"73747573", x"706D6C6C", x"6B69696A", x"69686869",
									 -- x"6F747B80", x"81807F7E", x"7B7B7C7D", x"80848B91", x"99999C99", x"8F8E9392", x"999D9891", x"95A1A8AA",
									 -- x"B2B0B3B6", x"B6BBC0C1", x"C5C2C0C0", x"C8C7CBE4", x"FAF7F2F2", x"FAFFFFFF", x"FFF3DDD1", x"C2AA9380",
									 -- x"7C736D69", x"6563615C", x"5A575753", x"4C494744", x"47424449", x"4A4B4E4F", x"484E5557", x"56585E65",
									 -- x"66656461", x"5B565658", x"5657585A", x"5A5B5B5B", x"58595957", x"57575653", x"53525151", x"504D4B4A",
									 -- x"4C4B4A49", x"47464342", x"43444443", x"4241403E", x"3B393633", x"312F2C2B", x"27242221", x"201D1C1C",
									 -- x"1D1C1A18", x"16151414", x"16131111", x"1212110F", x"0F101010", x"0F0E0C0B", x"110F0D0D", x"0E0E0C0A",
									 -- x"0F0E0E0E", x"0E0E0E0D", x"0D0C0D0D", x"0E0D0E0E", x"0F0F1010", x"0F0E0E0E", x"0E0F100E", x"0C0C0D0F",
									 -- x"0B0C0D0F", x"10100F0E", x"0D0D0D0C", x"0C0C0C0C", x"0B0B0B0B", x"0B0C0D0E", x"0E0E0E0D", x"0D0C0C0B",
									 -- x"0B0C0D0E", x"0E0D0C0C", x"0C0D0D0D", x"0D0E0E0E", x"0C0C0C0C", x"0D0E0F10", x"100F0E0E", x"0E0F0F0F",
									 -- x"10101010", x"10101010", x"0F101112", x"12121213", x"12121112", x"12121313", x"15141414", x"14141312",
									 -- x"14141413", x"13131212", x"14141414", x"14131415", x"15151616", x"17171717", x"16161717", x"17171819",
									 -- x"1A1B1C1D", x"1D1E1F20", x"1E1F2021", x"21212223", x"23242526", x"27272626", x"2A2A2A2A", x"2A2A2B2B",
									 -- x"7F7D7B79", x"77777878", x"79797978", x"78797B7C", x"81808081", x"83848485", x"8182817F", x"7E7E7C79",
									 -- x"76736F6C", x"6A676463", x"5856524F", x"4D4D5052", x"51525455", x"56585B5C", x"5D5E6163", x"64646565",
									 -- x"68696B6E", x"72777A7B", x"7D7E7E7E", x"80838484", x"82868989", x"898A8B8C", x"8D919191", x"93918E8F",
									 -- x"9396999A", x"9A9A9997", x"9A99999A", x"9C9D9D9D", x"9DA09E97", x"9596948F", x"9392908D", x"8A878482",
									 -- x"81808082", x"83858483", x"8687898B", x"89858588", x"85848383", x"817E7E7F", x"7F7F8185", x"84817E7D",
									 -- x"77767576", x"78787776", x"7A767471", x"6B6A6C6A", x"66666166", x"68656967", x"67666362", x"61616263",
									 -- x"61605E5B", x"5B5C5E5D", x"59585858", x"58595959", x"57595958", x"5656595C", x"5B5C5C5B", x"59595A5B",
									 -- x"5E5E5E5D", x"5D5D5F60", x"66686B6D", x"70737779", x"7E7F7E7C", x"77747271", x"6E6E7072", x"716F6E6E",
									 -- x"71778086", x"88868482", x"7B818586", x"8A939999", x"96999E9B", x"90909898", x"A7A6A09E", x"A5AEB9C6",
									 -- x"C1BEBFC1", x"C3C8CDCC", x"CBCED0CC", x"CECED7F3", x"FFFFFDFB", x"FEFEFDFE", x"FDF4DFD0", x"C3B09A83",
									 -- x"7D76716B", x"63605E59", x"58545350", x"4A484846", x"48485159", x"58565759", x"51545757", x"56575A5D",
									 -- x"5F5F5E5C", x"58535152", x"51515151", x"52535353", x"53545453", x"5252504D", x"4E4E4D4C", x"4B4A4846",
									 -- x"47464543", x"42413F3E", x"40404141", x"3F3D3B39", x"35333230", x"2F2D2B2A", x"27252322", x"211E1D1D",
									 -- x"1C1B1A19", x"17151312", x"14120F0F", x"1112110F", x"11100F0E", x"0E0D0D0D", x"0E0C0B0C", x"0E100F0E",
									 -- x"0E0D0D0D", x"0D0E0D0D", x"0C0D0D0C", x"0C0C0C0C", x"0F0E0C0C", x"0D0E0D0C", x"0D0E0E0C", x"0A0A0D10",
									 -- x"0B0B0B0C", x"0E0E0E0D", x"0D0D0D0C", x"0B0B0A0A", x"0B0B0B0B", x"0A0B0C0D", x"0A0B0C0C", x"0C0B0A0A",
									 -- x"0B0B0C0D", x"0D0D0C0C", x"0D0C0D0D", x"0D0D0D0E", x"0B0B0C0D", x"0E0E0D0D", x"0F0E0E0E", x"0F0F0E0E",
									 -- x"0E0D0D0E", x"0E0E0F10", x"0F0F1011", x"13131312", x"10111112", x"12111110", x"13121212", x"13131211",
									 -- x"10101112", x"13141515", x"13131413", x"13141617", x"17171818", x"18181818", x"16161718", x"1818191A",
									 -- x"191A1B1C", x"1C1D1E1F", x"20212121", x"21222324", x"24252626", x"27272828", x"2C2B2928", x"28292A2A",
									 -- x"7F7D7B78", x"76767778", x"77767473", x"73747473", x"76757577", x"797A7B7C", x"7C7D7C7A", x"7B7E7C78",
									 -- x"7472706F", x"6B666362", x"5955514E", x"4C4B4D4F", x"4E505151", x"52555859", x"595A5C5F", x"605F6061",
									 -- x"65666869", x"6D717272", x"76777776", x"787C7F7F", x"7C7E8081", x"81828485", x"84898A89", x"8C8C8A8B",
									 -- x"8D909291", x"90919292", x"94949291", x"93959594", x"94959491", x"8F908E8A", x"8B8A8986", x"827F7E7E",
									 -- x"7C7B7A7B", x"7D7E7E7D", x"7A7D8387", x"86828285", x"8684807D", x"7976787B", x"7B7A7C80", x"807B7776",
									 -- x"73737477", x"7A7A7774", x"74727474", x"706F6E6A", x"6C696469", x"6C6A6D6C", x"69696969", x"69686767",
									 -- x"6463615D", x"5C5D5E5D", x"5A595755", x"55545453", x"54545451", x"4F505356", x"54585958", x"56575B5E",
									 -- x"5B5C5E5E", x"5E606264", x"6B6F7478", x"7A7D8184", x"88888785", x"837F7C7A", x"74747578", x"79787676",
									 -- x"787B8086", x"898B8D8D", x"89909492", x"979FA19C", x"95999E9D", x"9A9DA4A7", x"B4B1AEB3", x"B9B7C5E3",
									 -- x"D4CECCD0", x"D5DCDFDB", x"D8D4D2D2", x"D8DCE0F3", x"EFFAFFFE", x"FEFDFCFF", x"FFF7E0D0", x"BEA89B8F",
									 -- x"847E786F", x"65615F5A", x"5752504F", x"4B4A4B4A", x"4C505E68", x"655E5D5E", x"5C5A5754", x"5457595A",
									 -- x"57565757", x"544F4C4B", x"4D4C4C4C", x"4D4D4D4D", x"4F50504E", x"4E4E4C4A", x"4A4A4745", x"44454443",
									 -- x"42413F3E", x"3E3E3D3D", x"3D3C3C3D", x"3C383535", x"32323130", x"302E2C2B", x"28252323", x"211F1D1D",
									 -- x"19181817", x"17151312", x"12110F0F", x"1010100F", x"100F0E0D", x"0D0D0E0E", x"0E0D0C0C", x"0E0F0E0E",
									 -- x"0D0D0C0C", x"0C0D0D0C", x"0C0D0D0C", x"0B0C0C0B", x"0F0D0B0B", x"0D0F0D0C", x"0C0C0C0B", x"0A0A0C0E",
									 -- x"0C0C0B0C", x"0C0C0C0B", x"0C0C0C0C", x"0A090909", x"0B0B0B0B", x"0A0A0B0C", x"0A0B0C0D", x"0D0C0B0A",
									 -- x"0D0C0B0A", x"0A0C0D0E", x"0D0C0C0D", x"0D0C0C0D", x"0D0D0E0F", x"0E0D0C0B", x"0E0E0E0E", x"0F0F0E0D",
									 -- x"0D0C0C0D", x"0E0F1113", x"10101012", x"13131210", x"11111313", x"13121110", x"12121213", x"13131312",
									 -- x"10101112", x"13141415", x"13151515", x"15171919", x"17171717", x"16161617", x"17181919", x"19191A1B",
									 -- x"1B1B1C1D", x"1D1D1E1F", x"1F202120", x"21232525", x"23242627", x"27292A2B", x"2C2B2B2A", x"2B2A2928",
									 -- x"7D7C7B7B", x"7B7A7775", x"76757371", x"73757370", x"716F7073", x"74747475", x"7777787A", x"7A797776",
									 -- x"74727172", x"70696361", x"5C585553", x"524F4F50", x"4E505252", x"53555757", x"5757585A", x"5B5A5C5F",
									 -- x"61636465", x"676A6C6B", x"6D6F7170", x"7275797A", x"7979797A", x"7B7D7E7F", x"7D828281", x"84858586",
									 -- x"85888A88", x"87898B8C", x"8D8D8B8A", x"8B8D8C8A", x"8B8A8A89", x"8A898886", x"8382817E", x"7A787778",
									 -- x"75737273", x"76787979", x"777A8188", x"88838183", x"83817E7C", x"78757578", x"7776787B", x"78737172",
									 -- x"71727376", x"797A7B7A", x"73717576", x"73716F6B", x"6F6C676D", x"6F6D7273", x"71727374", x"73727170",
									 -- x"6B6B6A67", x"65656463", x"5F5D5957", x"56555352", x"54535250", x"50505254", x"53575958", x"585C6062",
									 -- x"60616363", x"64676B6E", x"74797F83", x"8485888A", x"8E8D8D8D", x"8C898581", x"817E7D7F", x"81828181",
									 -- x"81828487", x"8C92989B", x"9B9F9F9E", x"A1A5A49F", x"9CA2A5A9", x"AFB3B4B5", x"BBBDBBC0", x"C6C3CEE9",
									 -- x"EAE6E5E4", x"E1E2E4E2", x"E4D7D3D4", x"D8D7D7E1", x"E7F2F7F6", x"F8F9F9FA", x"FBF2DECF", x"BEAAA29B",
									 -- x"91897F74", x"6A66645E", x"5A545252", x"4F4F504F", x"53586772", x"6C625F5F", x"5F5C5752", x"53555654",
									 -- x"504F5050", x"4F4B4847", x"4A494848", x"48494948", x"494A4A48", x"48494846", x"44444340", x"3F40403D",
									 -- x"3C3B3A3A", x"3B3B3A3A", x"38373738", x"37343233", x"32323131", x"302E2B2A", x"28252322", x"211E1D1D",
									 -- x"19181616", x"16151412", x"12111010", x"0F0F0F0F", x"0E0E0D0C", x"0C0D0E0F", x"0F0F0E0D", x"0C0C0B0B",
									 -- x"0D0C0B0B", x"0C0C0C0C", x"0B0D0D0B", x"0B0C0C0B", x"0D0C0C0D", x"0E0E0D0C", x"0C0C0B0B", x"0B0A0A0B",
									 -- x"0D0C0C0C", x"0D0C0B0A", x"0A0B0C0C", x"0A090909", x"090A0B0B", x"0B0B0B0B", x"0C0C0D0D", x"0D0C0C0B",
									 -- x"0D0C0B0A", x"0A0C0D0E", x"0D0C0B0D", x"0D0B0B0D", x"0D0E0E0E", x"0E0D0C0C", x"0E0E0D0D", x"0E0E0E0D",
									 -- x"0F0D0C0E", x"0E0F1114", x"10111313", x"13121111", x"12121313", x"13121110", x"12121314", x"14141312",
									 -- x"13131313", x"12121111", x"0E111110", x"11131514", x"15161514", x"13121314", x"16161718", x"18191A1B",
									 -- x"1B1C1E1E", x"1F1F2020", x"1E212222", x"22242424", x"24252728", x"28292A2C", x"2B2B2B2C", x"2E2E2C2B",
									 -- x"7F7B7777", x"78797774", x"73727070", x"7376746F", x"716F7174", x"75737273", x"7371747A", x"7A737175",
									 -- x"75727275", x"746E6661", x"615E5C5C", x"5A575555", x"54575755", x"54545452", x"55535355", x"5555585C",
									 -- x"5A5D5F60", x"62666766", x"696B6D6B", x"6B6D6E6F", x"76747374", x"7677797A", x"787C7B79", x"7C7E7E80",
									 -- x"7C7F8282", x"81828384", x"84848483", x"84868481", x"89858383", x"82807E7E", x"7E7D7A77", x"74727171",
									 -- x"6E6D6C6E", x"71747677", x"7E7F858E", x"908A8685", x"8080817F", x"7B757374", x"7676797A", x"76707075",
									 -- x"71727375", x"777B7F82", x"7C767270", x"6C6F7373", x"6D6C696F", x"716F7679", x"7A7A7B7B", x"7A7A7979",
									 -- x"74757470", x"6D6B6865", x"63615D5B", x"59585655", x"55555453", x"53545556", x"56595A5A", x"5C616566",
									 -- x"68696A6A", x"6B6F7478", x"888D9396", x"96949597", x"9A9A9A9B", x"9C99938D", x"908B8687", x"898B8B8C",
									 -- x"8A89898B", x"90989FA4", x"A3A1A1A3", x"A6A8A7A5", x"A8AFB2B9", x"C7C9C1BE", x"BFCAC7C4", x"CED4D8E4",
									 -- x"E6EAF0EE", x"E6E5EDF3", x"F0E5E8E5", x"D7CBCDDE", x"E3E7E3DF", x"E3E6E4E1", x"E7E5D6CB", x"C1B8B0A2",
									 -- x"998E8275", x"6C6A6760", x"5E575556", x"54545453", x"595D6B76", x"70645F5E", x"5C5A5550", x"50504E4A",
									 -- x"4D4B4B4B", x"4A474545", x"46444343", x"44444443", x"44454443", x"43454442", x"3E40403F", x"3E3E3B37",
									 -- x"38383737", x"38373635", x"35333334", x"33313133", x"30302F2E", x"2D2A2725", x"27252222", x"211E1C1D",
									 -- x"1B191716", x"15151413", x"13131211", x"0F0E0F10", x"0C0C0C0C", x"0D0D0E0E", x"0C0D0D0C", x"0C0C0C0D",
									 -- x"0D0C0B0B", x"0B0C0C0C", x"0A0C0C0B", x"0B0D0D0B", x"080A0C0C", x"0C0B0A0A", x"0B0B0B0B", x"0C0B0907",
									 -- x"0B0C0C0D", x"0E0E0C0B", x"090A0C0C", x"0A09090A", x"08090A0B", x"0B0B0B0B", x"0B0B0B0B", x"0A0A0A0A",
									 -- x"0B0B0C0C", x"0D0D0C0C", x"0D0B0B0D", x"0C0B0A0C", x"0B0B0C0C", x"0C0D0D0D", x"0F0E0C0C", x"0D0D0E0E",
									 -- x"110D0C0C", x"0C0C0E11", x"0E111414", x"12111113", x"13131312", x"12111111", x"10101113", x"1312110F",
									 -- x"13131313", x"13121111", x"10131312", x"12151615", x"16161614", x"12111214", x"12131416", x"17181A1B",
									 -- x"191B1D1E", x"1F202122", x"20232524", x"23242422", x"25262829", x"2929292A", x"2B2A2A2C", x"2F313131",
									 -- x"7E7D7B78", x"75757779", x"72707675", x"72706D71", x"71717271", x"71717173", x"70757A79", x"74727478",
									 -- x"72727374", x"73706D6A", x"65646466", x"64616061", x"5F5C5C5B", x"58565450", x"52505052", x"51505359",
									 -- x"5355595D", x"5C5B5F64", x"66636367", x"6865686E", x"6A6D6D6C", x"6D71716E", x"6F707375", x"75737579",
									 -- x"7879797B", x"7D7C7B79", x"7D7D7E7E", x"7E7E7E7E", x"7A7A797A", x"7A787573", x"76777672", x"706E6D6B",
									 -- x"6D6B6968", x"6A6E7376", x"7E858890", x"928E8F8A", x"898A8782", x"7F807D78", x"78777778", x"76757576",
									 -- x"72747576", x"7A7F807F", x"78777674", x"716E7074", x"76737070", x"72777E82", x"81808082", x"8484827F",
									 -- x"7C807F77", x"74746D63", x"615F5E5C", x"5B585757", x"54595854", x"585C5A58", x"5C616161", x"65696C70",
									 -- x"72737579", x"7B7F868D", x"97A6ADAB", x"ABAAA5A0", x"A5AAADAA", x"A49E9D9E", x"9C989595", x"94939393",
									 -- x"8E8A8C92", x"979FA7AA", x"ACAEA8A6", x"ACAEB2BE", x"BDC4C4C1", x"C8D3CEBF", x"C7CFD1D3", x"D8DAE0ED",
									 -- x"E7E9F3F7", x"F2F3F8F8", x"F8EFF4FA", x"EBD8D3D5", x"DADBD8D1", x"D2DEE2DA", x"D4CFCDCB", x"C3BBB1A8",
									 -- x"9C918880", x"76706D6A", x"675E5A5A", x"58595956", x"5F686E6B", x"645F5B57", x"5E59534E", x"4E4F4C46",
									 -- x"48474646", x"48474440", x"42403E3E", x"3F403F3E", x"40403F3E", x"3D3D3D3D", x"3D3C3B3A", x"39383635",
									 -- x"35323131", x"3232302F", x"31313130", x"302F2F2F", x"2C2D2D2C", x"2A282726", x"2121201F", x"1F1E1C1A",
									 -- x"1C191514", x"16161512", x"12111010", x"0E0C0D0E", x"0F0D0C0B", x"0B0C0D0D", x"0E0D0B0A", x"0A0B0C0D",
									 -- x"0F0E0C0B", x"0C0C0C0B", x"0B0A0A0B", x"0C0C0A08", x"0D0C0B0A", x"0A0B0B0C", x"0B0B0A08", x"08080A0B",
									 -- x"0A0A0A0A", x"0A0A0B0C", x"0D0C0A0A", x"0B0B0907", x"0808090A", x"0B0B0B0B", x"090A0A0B", x"0B0B0A0A",
									 -- x"0B0B0C0B", x"0A090A0B", x"0C0C0C0C", x"0C0B0A09", x"0C0B0B0D", x"0E0E0C0A", x"0D0D0D0D", x"0D0D0E0E",
									 -- x"110F0D0C", x"0C0D0D0E", x"11100E0E", x"0F111213", x"16121011", x"12111010", x"0E101212", x"11111213",
									 -- x"11100F10", x"13131211", x"12131314", x"13131415", x"16151413", x"14141514", x"18181818", x"1718191A",
									 -- x"18191A1A", x"1B1C1F21", x"20212225", x"25222121", x"23272A29", x"27272A2E", x"2D2D2E30", x"2F2D2F32",
									 -- x"7A7B7C7B", x"79787777", x"72707574", x"74757378", x"75726F6F", x"72737271", x"70737677", x"75747576",
									 -- x"7777797A", x"7A787573", x"6D6E7072", x"706B6766", x"67626261", x"5E5C5953", x"53515050", x"504E4E4F",
									 -- x"4B4B4F53", x"5555585B", x"5C5D5D5F", x"60626466", x"6868686A", x"6B6A6A6A", x"6A696A6C", x"6D6C6D6F",
									 -- x"70707173", x"75757573", x"73757677", x"76777879", x"75747374", x"7473716F", x"6F70706D", x"6B6C6E6E",
									 -- x"6E6D6A69", x"6A6D7174", x"7D838690", x"96979996", x"9697948D", x"89898987", x"82818182", x"817F7F81",
									 -- x"84858685", x"86898B8A", x"8085857E", x"76747576", x"7A7A7E84", x"88898B8D", x"89898A8A", x"89888686",
									 -- x"86827D7A", x"756E6968", x"64646361", x"5F5D5B5A", x"5C62615E", x"60616061", x"63696C6F", x"767C7E82",
									 -- x"80818488", x"8C919AA2", x"ACB7BCBA", x"BCBDBAB8", x"B7B7B7B7", x"B8B7B4B1", x"ADB0ACA3", x"A0A39F96",
									 -- x"99989BA0", x"A4ACB3B3", x"BABBB6B7", x"BEC1C3CB", x"CECFCDCB", x"CDD2D1CD", x"CFD8E0E4", x"E5E2DFE1",
									 -- x"E0DBE3F1", x"F7F5F6F8", x"F4F4FAFA", x"EDDFD9D8", x"DEDDDDDA", x"D7DBE1E0", x"E0DBD6D1", x"C9C3BDB4",
									 -- x"A3978D86", x"7D797874", x"6E666160", x"5E5D5D5B", x"61696D69", x"625E5956", x"55534F4A", x"494A4846",
									 -- x"47454343", x"4443413E", x"3D3B3A3A", x"3C3C3C3B", x"3E3D3B3A", x"3A3A3B3C", x"39383737", x"36353332",
									 -- x"322F2D2D", x"2E2E2D2C", x"2D2D2D2D", x"2D2D2D2C", x"2A2A2928", x"26252423", x"20201F1F", x"1E1D1B1A",
									 -- x"1A171413", x"14141210", x"100E0D0D", x"0C0A0A0C", x"0D0C0C0C", x"0C0D0D0D", x"0D0D0C0B", x"0B0B0B0B",
									 -- x"0C0B0B0B", x"0C0C0C0B", x"0D0C0C0D", x"0E0D0C0A", x"0C0B0B0B", x"0A0B0B0B", x"0C0B0B0A", x"09090B0C",
									 -- x"0B0C0C0C", x"0B0B0C0D", x"0D0B0A0A", x"0B0B0A08", x"0B0B0B0B", x"0A0A0909", x"0808090A", x"0A0B0B0A",
									 -- x"0A0B0B0A", x"0A090A0B", x"0C0C0C0C", x"0C0B0B0B", x"0B0C0D0D", x"0C0C0B0B", x"0C0D0D0D", x"0D0E0F0F",
									 -- x"0F0E0D0C", x"0D0E0F0F", x"11101010", x"12131313", x"110E0D0E", x"10100F0F", x"0F0F1011", x"12121111",
									 -- x"11101011", x"12121211", x"13131414", x"14151516", x"17151413", x"14151516", x"16161717", x"1819191A",
									 -- x"1A1A1B1B", x"1C1D2022", x"20212323", x"211F2023", x"26292B2A", x"28282A2D", x"2B2B2C2F", x"302F3032",
									 -- x"7D7C7A79", x"78777777", x"74717574", x"7679787C", x"7B787574", x"76787878", x"7B7B7C7D", x"7E7E7D7D",
									 -- x"7B7C7E80", x"81807E7D", x"7C7B7978", x"76727070", x"6C676665", x"615E5A53", x"5353514F", x"4F4E4B47",
									 -- x"4746484C", x"4F515152", x"51545656", x"575C5E5E", x"625F6065", x"66626264", x"66646465", x"67676768",
									 -- x"6768686A", x"6B6C6C6C", x"6B6E7070", x"70707274", x"72706F6E", x"6F6F6E6D", x"6B6D6C6A", x"696C7073",
									 -- x"71706F6D", x"6D6E7173", x"7E82848E", x"95989D9A", x"9B9E9D98", x"93939493", x"908F8F8F", x"8E8C8C8E",
									 -- x"9293918E", x"8C8D8F8F", x"858B8C85", x"8182827F", x"81838A92", x"94908D8F", x"8D8B8B8E", x"9192908E",
									 -- x"8D857C76", x"6F69686B", x"67676766", x"64636160", x"60656566", x"6A6B6C70", x"737A7F83", x"8B909396",
									 -- x"96969799", x"9CA1AAB1", x"B8BDBEBE", x"C1C2C1C3", x"C6C4C2C3", x"C6C6C4C1", x"BEC1BDB5", x"B3B5B0A5",
									 -- x"A9AAADB0", x"B3BABFBC", x"C1C2C1C6", x"CED1D2D6", x"DEDAD8D8", x"D6D4D6DA", x"DBE2EDF1", x"EEE7DDD1",
									 -- x"D4D7DEED", x"F8F8F6F9", x"F1F6F3E8", x"E0DDDCDD", x"E0E1E9EE", x"E7E0DEDF", x"DFDCD8D1", x"C8C4BFB7",
									 -- x"A79C938F", x"8986837F", x"776E6866", x"6261615E", x"666B6E69", x"625D5853", x"51514F4A", x"47464646",
									 -- x"4543403F", x"3F3E3C3A", x"39373637", x"38393837", x"3B393736", x"35363738", x"33333232", x"3231302E",
									 -- x"2D2B2929", x"2A2B2B2A", x"2C2C2B2B", x"2B2A2A2A", x"26262523", x"22212020", x"1F1E1D1D", x"1D1B1A18",
									 -- x"18151211", x"1211100E", x"0F0E0D0D", x"0C0A0A0B", x"0A0B0C0D", x"0D0D0D0C", x"0D0D0C0C", x"0B0A0A09",
									 -- x"09090A0B", x"0C0C0B0A", x"0C0B0B0B", x"0C0B0A09", x"0A0B0B0B", x"0B0B0B0B", x"0C0C0C0B", x"0B0A0B0C",
									 -- x"0B0C0C0C", x"0C0C0C0D", x"0C0B0A0B", x"0B0B0A09", x"0C0C0B0A", x"0A090909", x"07080809", x"090A0A0A",
									 -- x"090A0A0A", x"0A0A0B0C", x"0C0C0C0B", x"0B0C0C0C", x"0B0C0E0D", x"0B0A0B0C", x"0C0D0E0E", x"0E0F1011",
									 -- x"0E0E0D0E", x"0F101010", x"11111213", x"14141413", x"100D0C0E", x"10101010", x"100F0F10", x"1212100E",
									 -- x"10111212", x"12111112", x"14131314", x"16171717", x"17161414", x"14151617", x"16161618", x"1A1B1B1A",
									 -- x"1B1B1C1C", x"1D1E2123", x"20212222", x"1F1D2025", x"28292A2A", x"29292B2C", x"2D2D2E2F", x"2F2E2D2E",
									 -- x"7F7E7C7B", x"7A797777", x"78757877", x"787C797C", x"7B7E7F7D", x"7A7A7E83", x"80808081", x"82828180",
									 -- x"81828385", x"86868584", x"8683807E", x"7C7A7878", x"726F6E6C", x"65615C56", x"5455534E", x"4D4E4D48",
									 -- x"4A494A4C", x"4F4F4E4E", x"4C4E5051", x"52555758", x"5957595C", x"5E5D5C5E", x"61606061", x"62626364",
									 -- x"63636363", x"64646565", x"67696B6B", x"6A6A6D6F", x"706D6B69", x"6A6A6A69", x"6A6C6B69", x"686B6F72",
									 -- x"71717170", x"6F6F7172", x"7E83838A", x"8F909594", x"94989A99", x"97969594", x"94939393", x"92909092",
									 -- x"99989691", x"8D8C8E90", x"87888887", x"898C8984", x"8A8A8E91", x"8D848286", x"8A85858E", x"9AA09C94",
									 -- x"8E897D6F", x"686A6D6D", x"6C6D6D6C", x"6B6B6B69", x"6A6C6C70", x"77797B81", x"89919697", x"9B9EA0A5",
									 -- x"A7A6A5A5", x"A7ADB5BB", x"C3C4C3C5", x"C8C7C5C8", x"CECFCECD", x"CCCBCACA", x"CDCAC9CA", x"CAC6C0BC",
									 -- x"BABBBEBF", x"BFC6C9C5", x"C6C8CCD3", x"DBDDDEE1", x"E6E3E3E5", x"E3DEDFE5", x"E4E8F2F5", x"F1EEE3D1",
									 -- x"D0E2EBED", x"F5FAFAFB", x"F9FDF2E5", x"E3E5E5E9", x"E7E7EFF5", x"EEE4DDD9", x"D1D3D3CD", x"C2BFBCB6",
									 -- x"AEA49E9B", x"97938E87", x"7D746F6C", x"67656461", x"696D6E69", x"635E5852", x"52514F4B", x"46444343",
									 -- x"413F3D3C", x"3B3B3937", x"37363535", x"36363535", x"38363533", x"32313232", x"2E2E2E2E", x"2E2E2D2C",
									 -- x"29292929", x"2A2C2C2A", x"2A2A2928", x"27262525", x"2322201F", x"1E1E1E1D", x"1C1C1B1B", x"1B1A1817",
									 -- x"16141211", x"10100E0D", x"0F0D0C0D", x"0D0B0A0B", x"0A0B0C0D", x"0D0C0C0C", x"0C0C0C0B", x"0B0A0A09",
									 -- x"0808090A", x"0B0B0A09", x"0A090909", x"09090808", x"0A0A0B0C", x"0C0C0B0B", x"0B0C0C0C", x"0B0B0B0B",
									 -- x"0A0B0C0C", x"0B0B0C0C", x"0B0B0A0B", x"0B0B0A09", x"0B0A0A09", x"090A0A0B", x"09090909", x"09090808",
									 -- x"0A0A0A0A", x"0B0B0C0D", x"0D0C0B0B", x"0B0C0D0E", x"0C0C0D0C", x"0B0B0D0E", x"0D0E0F0F", x"0F101011",
									 -- x"0F0F0F0F", x"1010100F", x"12121213", x"14141312", x"100E0E0F", x"10100F10", x"10101011", x"1212100F",
									 -- x"0F111313", x"11111213", x"13131314", x"16171717", x"19171514", x"15161717", x"18171719", x"1C1D1C1B",
									 -- x"1B1B1C1C", x"1E202224", x"20212223", x"211F2123", x"26262728", x"292B2C2D", x"2F2F2F2F", x"2F2E2E2D",
									 -- x"7F808282", x"817F7C7A", x"7D7B7F7D", x"7D807C7C", x"7A7E8180", x"7D7D8084", x"81828384", x"84858586",
									 -- x"8888898A", x"8B8B8A89", x"87888A8A", x"8985807B", x"7C7A7A77", x"6E68645F", x"5657544E", x"4B4D4E4D",
									 -- x"4C4C4D4E", x"4E4E4D4C", x"4C4A4B4F", x"504E4F53", x"51535454", x"56585855", x"57595A5A", x"595A5C5E",
									 -- x"5E5E5E5E", x"5E5F6061", x"62646564", x"63636567", x"6A676564", x"64656665", x"66686866", x"66686B6D",
									 -- x"6D6E6F6E", x"6D6D6F71", x"7A818388", x"89888E8F", x"8D8F9192", x"9293918E", x"8D8D8D8F", x"8F8D8E90",
									 -- x"9493918C", x"8886888B", x"8A87878A", x"8A868383", x"8B8B8C8B", x"82797A80", x"8582858F", x"9CA29E97",
									 -- x"8F887A6C", x"676B7175", x"76777775", x"75777776", x"7B7C7B7E", x"868A8B90", x"9CA5A8A7", x"A7A7AAB0",
									 -- x"B0B0B0B1", x"B4BBC3C8", x"CCCECFD3", x"D7D4D0D2", x"D6D6D7D7", x"D7D6D6D6", x"D9D9DDE2", x"E3DCD3CD",
									 -- x"C9C9CCCC", x"CBD1D5D2", x"D5D7DFE6", x"E9EAECEE", x"EDECEDEE", x"EDEBEBEC", x"EAECF4F7", x"F6F7F0E0",
									 -- x"DAECF3F2", x"F6FAFAFD", x"FCFEF8F4", x"F7F5EDEB", x"F0ECEBEA", x"E6E3DDD5", x"CACDD0CB", x"C2BFC0BC",
									 -- x"BCB1ABA8", x"A29D9790", x"837B7672", x"6C696865", x"686B6C69", x"65615A54", x"524F4C49", x"4643403E",
									 -- x"3D3C3B3A", x"3A383635", x"35343433", x"33333231", x"32323130", x"2F2E2D2D", x"2B2B2B2C", x"2C2C2B2A",
									 -- x"28292A29", x"292B2A27", x"25252423", x"22212020", x"201F1E1D", x"1D1D1D1C", x"1A191919", x"19181615",
									 -- x"14141211", x"100F0E0E", x"0E0B0B0C", x"0C0A0909", x"0B0C0D0D", x"0C0C0C0C", x"0C0C0B0A", x"0A0A0B0B",
									 -- x"09090909", x"0909090A", x"0A0B0B0B", x"0A0A0A0A", x"0A0B0C0D", x"0D0D0C0B", x"0A0B0C0C", x"0B0A0A0A",
									 -- x"090A0B0C", x"0C0C0C0D", x"0B0B0B0B", x"0B0B0A09", x"09090808", x"09090A0A", x"09090909", x"09090909",
									 -- x"0A0A0A0B", x"0B0C0D0D", x"0D0C0B0B", x"0B0C0E0E", x"0D0C0B0B", x"0D0E0E0E", x"0D0E1010", x"10101011",
									 -- x"0F0F0F10", x"11111010", x"12121111", x"11111111", x"0E0D0D0F", x"100F0F10", x"10121313", x"12111111",
									 -- x"0F111313", x"11111214", x"15141414", x"15151515", x"19181615", x"15161617", x"1A19181A", x"1C1D1C1A",
									 -- x"1B1B1B1D", x"1F212324", x"20202124", x"25232222", x"24242526", x"282A2B2C", x"2C2D2E2E", x"30313333",
									 -- x"84858685", x"8586888A", x"87878B87", x"86888282", x"81808182", x"84858381", x"81838687", x"87888A8C",
									 -- x"8C8C8C8D", x"8E8E8E8D", x"8D8E8E8E", x"8E8D8884", x"8280807C", x"736E6A66", x"5C5C5852", x"4D4D4F50",
									 -- x"4B4D4E4E", x"4E4E4D4B", x"4E4A4A4E", x"4E4A4A50", x"4E51514E", x"4F53524E", x"4F525453", x"51525556",
									 -- x"56575859", x"595A5C5D", x"5F5F5F5E", x"5E5E5F60", x"64626060", x"61636362", x"61636464", x"64676868",
									 -- x"686A6C6C", x"6B6B6D70", x"717A7F85", x"85858C8E", x"8B8A8A8A", x"8B8C8C8B", x"8686888A", x"8B8B8C8E",
									 -- x"8E8C8A88", x"86848588", x"8786888A", x"857D7D83", x"82838583", x"7E797A7F", x"7F838A90", x"94959493",
									 -- x"9180716D", x"6A686F7A", x"7F81817F", x"7F818280", x"8486878A", x"9297999C", x"A4ADB2B0", x"AFAEB0B6",
									 -- x"B7B8B9BA", x"BEC5CBCE", x"CFD4D8DE", x"E4E2DDDE", x"DBD8D6DA", x"E0E4E3E1", x"DBE6EFF0", x"F2F2E8DB",
									 -- x"D5D3D5D7", x"D6DADFDF", x"E5E5EDF3", x"F1F1F4F3", x"F2F2F2F1", x"F0F1F1F1", x"F2F4F8FA", x"FAF9F3E9",
									 -- x"EBEBEEF5", x"FBF9F8FE", x"FEFCFAFC", x"FFFDF2EB", x"EDEAE8E5", x"E4E5DFD3", x"CBC9CAC8", x"C3C3C5C4",
									 -- x"C7BCB4AE", x"A7A29D97", x"89817D79", x"736E6C69", x"676A6A67", x"66635D56", x"514D4948", x"4744403D",
									 -- x"3B3A3A39", x"38363533", x"31313130", x"2F2E2D2D", x"2C2C2D2D", x"2D2C2B2B", x"2929292A", x"2A2A2928",
									 -- x"27292927", x"25262522", x"21212020", x"201F1F1F", x"1F1D1C1C", x"1C1C1B1A", x"18171717", x"17161514",
									 -- x"12121211", x"0F0E0E0E", x"0E0C0B0C", x"0D0B0A09", x"0B0D0E0E", x"0C0B0C0C", x"0C0C0B0A", x"0A0B0B0C",
									 -- x"0B0A0A08", x"0708090B", x"0A0B0B0B", x"0B0A0B0C", x"0A0B0C0C", x"0D0C0B0B", x"0A0B0B0B", x"0A0A0A0A",
									 -- x"0A0B0C0D", x"0D0C0D0D", x"0C0C0C0B", x"0B0A0909", x"09090908", x"08080808", x"08080808", x"08090A0A",
									 -- x"0B0A0A0A", x"0C0C0D0C", x"0D0C0B0B", x"0B0C0D0E", x"0E0C0B0B", x"0D0F0E0D", x"0D0F1010", x"10101010",
									 -- x"0E0E0E10", x"11121211", x"1311100F", x"10101111", x"0E0D0E11", x"11111113", x"11121313", x"11101113",
									 -- x"10121313", x"12111214", x"16161615", x"13121213", x"19181616", x"16161616", x"19191819", x"1A1B1A19",
									 -- x"1B1B1C1E", x"21232324", x"21202125", x"27262423", x"24242526", x"2728292A", x"2B2E302F", x"30313334",
									 -- x"8D909292", x"9192979B", x"96969A95", x"91918C8C", x"8C8A898A", x"8C8B8884", x"81828486", x"8687898B",
									 -- x"8E8E8E8F", x"90919191", x"9393918F", x"8F91908D", x"8681807E", x"7875716B", x"67635F5B", x"57545355",
									 -- x"51525252", x"5455534E", x"504E4D4E", x"4C4A4B4E", x"4E4D4C4C", x"4C4D4D4C", x"4C4F504F", x"4E4F5050",
									 -- x"51525354", x"55555758", x"5B5A5959", x"5A5C5C5C", x"605E5D5D", x"5E5E5D5C", x"5D5E5F5F", x"61646462",
									 -- x"60636566", x"6566696B", x"6870757C", x"7E7E8587", x"87868686", x"85858586", x"82828385", x"86858789",
									 -- x"8B898889", x"88878789", x"84828383", x"817D7D7F", x"7A7C7D7C", x"7C7D7E7D", x"7C838A8D", x"8C8B8C8E",
									 -- x"917E6F6D", x"6C696F7A", x"83878988", x"898C8C89", x"89919596", x"9CA1A3A6", x"A9B3B9BA", x"BAB8B6B7",
									 -- x"B9BBBDBE", x"C1C7CBCC", x"CFD8DFE5", x"ECECE9E9", x"E0DDDADB", x"E1E6E7E7", x"DEEAF2F3", x"F5F8F3E9",
									 -- x"E1DDE0E4", x"E2E2E7E9", x"ECE9EEF3", x"F0F1F3F0", x"F5F4F4F5", x"F4F2F3F5", x"F9FBFBFB", x"FCF8F3F1",
									 -- x"F4EBEDF7", x"FBFAFBFE", x"FFFFFDFF", x"FFFFFAF0", x"E2E4E8E8", x"E7E7E2D7", x"D0C7C6CA", x"CACAC9C7",
									 -- x"C8BFB9B5", x"ADA7A29D", x"938C8885", x"7D777470", x"6D6D6B67", x"66655F58", x"524E4A4A", x"4945413F",
									 -- x"3B3A3937", x"35343332", x"2E2E2E2E", x"2D2B2B2A", x"29292929", x"29292929", x"27272728", x"28282726",
									 -- x"26282722", x"2122221F", x"1F1F1F1F", x"1F1F1E1E", x"1E1C1B1A", x"1B1A1816", x"16161515", x"16151412",
									 -- x"0F101110", x"0E0D0D0E", x"0F0C0B0D", x"0E0C0A0A", x"0A0C0F0F", x"0E0C0C0D", x"0C0C0C0C", x"0B0B0B0B",
									 -- x"0B0B0A09", x"08080A0B", x"090A0A0A", x"0A0A0B0C", x"0A0B0B0B", x"0B0B0A0A", x"0A0B0B0B", x"0A0A0A0A",
									 -- x"0B0C0D0D", x"0C0B0B0B", x"0C0C0C0C", x"0A090908", x"0A0A0A09", x"09080807", x"08080707", x"08080909",
									 -- x"0B0A090A", x"0B0C0C0B", x"0C0C0B0B", x"0B0B0C0D", x"0D0C0C0C", x"0C0C0C0C", x"0C0E0F10", x"10101011",
									 -- x"0F0E0E0F", x"10111111", x"12111010", x"11111212", x"0F0F1013", x"13121214", x"11121111", x"11111212",
									 -- x"12131413", x"12111212", x"14151615", x"13121315", x"17161616", x"17171717", x"19191919", x"191A1A1A",
									 -- x"1C1D1E20", x"23242322", x"21202023", x"25252627", x"25262727", x"2727292A", x"2A2F3332", x"30303132",
									 -- x"9199A4A9", x"A7A3A1A1", x"A2A2A59E", x"98989292", x"92939391", x"8E8C8A8A", x"8A8A8B8B", x"8C8D8E8E",
									 -- x"90909192", x"94969797", x"94959695", x"9797948F", x"8D868382", x"807E7972", x"6F6A6665", x"625D5A5A",
									 -- x"5B5A5858", x"5C5E5A53", x"5152514D", x"4C4D4E4D", x"4D49484B", x"4C4A4A4D", x"4B4C4C4B", x"4C4E4D4A",
									 -- x"4F505252", x"52525354", x"56545354", x"575A5A59", x"5D5B5A59", x"59585654", x"59595959", x"5C5F5E5B",
									 -- x"585B5D5E", x"5D5E6164", x"636A6C73", x"75757B7B", x"7F818484", x"82808081", x"7F7E7F80", x"7F7E7E80",
									 -- x"817E7E80", x"817F7F80", x"85817C7B", x"7F817D76", x"7B7B7978", x"7C81807C", x"7E82888B", x"8B8B8D8E",
									 -- x"9386776E", x"6E717679", x"868B8F90", x"92969592", x"94A1A7A5", x"A7AAABAD", x"B0BAC0C3", x"C6C2BBB9",
									 -- x"B6B9BCBF", x"C3C9CCCC", x"CAD4DCE2", x"E9ECEAE9", x"E7E6E4E1", x"E0E2E7EC", x"E9EBEFF2", x"F3F2F2F4",
									 -- x"EDE8EAF0", x"EDEAEDF1", x"EEE8ECF1", x"EFF1F3EF", x"F6F5F8FC", x"FAF5F5FA", x"FAFDFAFA", x"FEFBF8FE",
									 -- x"F4EFF3F8", x"F8FCFFFE", x"FFFCFEFE", x"FCFFFAEB", x"DCDEE4E6", x"E3E3E4E0", x"D6C9C7D0", x"D4D3CDC7",
									 -- x"C5BFBEBD", x"B6AFA8A2", x"9E989490", x"88817E7A", x"75736E69", x"66655F58", x"524E4B4B", x"4844403F",
									 -- x"3C3B3835", x"33323232", x"2C2C2D2D", x"2C2A2A2A", x"29282726", x"26262627", x"26262626", x"26262524",
									 -- x"2426241F", x"1E212220", x"1E1D1D1D", x"1C1B1B1B", x"1D1B1A1A", x"1A191613", x"15151415", x"15141312",
									 -- x"0D0F100F", x"0D0C0C0D", x"0D0A090B", x"0C0B0908", x"080C0F11", x"0F0E0D0D", x"0C0D0D0D", x"0D0B0A09",
									 -- x"0A0B0B0A", x"09090A0C", x"090A0B0B", x"0A0B0C0E", x"0A0A0A0A", x"0A090909", x"0B0B0B0B", x"0A0A0A0B",
									 -- x"0A0B0C0C", x"0B090908", x"0C0D0D0C", x"0A090808", x"090A0A0A", x"0A090808", x"09080707", x"06070707",
									 -- x"0A090809", x"0A0B0A0A", x"0C0C0B0B", x"0B0B0B0C", x"0B0D0D0C", x"0A090A0B", x"0B0D0F10", x"11111111",
									 -- x"11100F0F", x"1010100F", x"11101011", x"12131313", x"100F1012", x"11101011", x"12110F0F", x"11121211",
									 -- x"14141413", x"12111110", x"10131615", x"13131518", x"15151516", x"17181817", x"1A1A1A1A", x"191A1B1C",
									 -- x"1E1E2022", x"24242321", x"22212021", x"2223272B", x"26272828", x"27282A2B", x"252D3232", x"30313233",
									 -- x"A8AEB4B6", x"B6B4B0AC", x"AFB1ADA5", x"A4A8A59D", x"9D9E9D9A", x"95929292", x"90909193", x"92908F8F",
									 -- x"91959694", x"959A9B9A", x"98979798", x"98969697", x"9091908C", x"88837E7A", x"7674706B", x"67656463",
									 -- x"65636162", x"6363605E", x"5C57524F", x"5051504E", x"4D4D4E4E", x"4D4D4D4E", x"4D4D4C4C", x"4B4B4A4A",
									 -- x"4C4F5150", x"4E4E5256", x"54535353", x"53525355", x"53555757", x"54535456", x"58575554", x"56595957",
									 -- x"57575554", x"55575B5E", x"59606468", x"6E716F70", x"71767A7B", x"79797A7A", x"7A797371", x"74757578",
									 -- x"787B7D7D", x"7A787878", x"75747679", x"77737478", x"7878747A", x"7D7B8183", x"7E818486", x"8484898F",
									 -- x"8F8C837C", x"7B7A7D85", x"89898E96", x"9C9F9E9E", x"A3ABAEAE", x"B2B5B4B4", x"B3BAC0C2", x"C1C1BEBC",
									 -- x"BEBAB9BD", x"C1C2C6CB", x"CFD4D7DA", x"E1E3E4E7", x"EAE9E8E6", x"E3E2E6EB", x"E6ECF1F2", x"F2F2F2F2",
									 -- x"F1F0EFF0", x"F2F3F2F1", x"F1F1F0EF", x"EFF1F4F6", x"F4F4F7FB", x"FCFAFAFC", x"FCFCFBFC", x"FDFDFBFA",
									 -- x"F5F7FBFD", x"FEFEFCFC", x"FFFCFDFF", x"FFFEF0DF", x"D4D3D8DD", x"DBDCDFE0", x"D9D0C9CB", x"D3D6D3CF",
									 -- x"C8C6C2BD", x"B8B2AEAC", x"A9A8A49D", x"97918A84", x"7F79746D", x"6765625A", x"56534E4A", x"4643403D",
									 -- x"3B3A3A38", x"3532302F", x"2C2A2C2C", x"28282928", x"25252424", x"23242627", x"22252625", x"25262421",
									 -- x"22222121", x"1F1E1C1B", x"1C1D1C1B", x"1A191A1A", x"1B191816", x"16151413", x"13141412", x"13151412",
									 -- x"110F0F0F", x"0E0C0C0D", x"0D0D0B0A", x"0A0B0C0C", x"0B0C0E0F", x"0E0D0D0E", x"0E0E0D0B", x"0A090A0B",
									 -- x"08090A0B", x"0B0B0A09", x"0B0A0A0A", x"0A0A0A0A", x"07080809", x"0A0A0A0A", x"0B0B0B0B", x"0C0C0A08",
									 -- x"090A0B0C", x"0B0A0908", x"080B0C0B", x"09080808", x"09080707", x"07070707", x"07090908", x"07080909",
									 -- x"090B0B0A", x"0B0C0C0A", x"0B09090A", x"0B0A0B0D", x"0D0C0B0A", x"0A0B0D0E", x"0C0D0F0F", x"0F0E0E0D",
									 -- x"0D0D0D0D", x"0E0E0E0E", x"0F101011", x"10100F0F", x"11111112", x"13131211", x"12100E10", x"13151412",
									 -- x"11131616", x"15131212", x"14131314", x"14151514", x"16161718", x"1919191A", x"191A1B1D", x"1D1D1D1C",
									 -- x"1A202424", x"23232220", x"22252122", x"23252B28", x"25272929", x"27262729", x"292B2A2D", x"31313238",
									 -- x"B4B9BDBF", x"BFBFBDBA", x"B9B7B5B3", x"B1B0AEAC", x"AEADABA7", x"A29D9998", x"97959596", x"97969596",
									 -- x"97989999", x"9DA09E98", x"9A999A9C", x"9D9A9898", x"93949492", x"908C857E", x"7B7A7773", x"716F6E6E",
									 -- x"6E6F6F6F", x"6C696664", x"615C5754", x"54545453", x"52525150", x"4F4E4E4F", x"4D4D4D4E", x"4E4E4E4D",
									 -- x"4A4C4E4D", x"4C4B4D4F", x"52504F50", x"4F4F5153", x"52504F50", x"53545351", x"5352504F", x"52555553",
									 -- x"53525150", x"50525456", x"585E5F61", x"66686768", x"6C707473", x"71707070", x"6E706F70", x"73716D6D",
									 -- x"71747676", x"74737375", x"75737376", x"76737377", x"76787577", x"79797E7B", x"797A7C7D", x"7E80878D",
									 -- x"8E8B8688", x"8D8D8889", x"8F91949A", x"A1A6A8A8", x"AEB3B4B4", x"B7B7B5B7", x"B4B8BBBC", x"BCBFC1C1",
									 -- x"BFBCBCC0", x"C2C3C6CA", x"CED5D8DB", x"DFE1E4EA", x"EDEBE9E8", x"E5E4E5E9", x"EBEEF1F2", x"F2F4F4F3",
									 -- x"EFF0F0F1", x"F2F2F3F3", x"F2F1F0F0", x"F1F3F4F5", x"F7F4F4F8", x"FCFDFDFE", x"FAF8F7F8", x"FBFBFAF9",
									 -- x"F9FBFDFF", x"FFFFFFFF", x"FFFBF9F9", x"F7F3E9DC", x"D1CCCDD1", x"D2D5D8D7", x"D7D0CACB", x"CED0CECD",
									 -- x"C5C5C3C0", x"BBB5B0AC", x"ACACA9A3", x"9C958E88", x"817A746E", x"67646159", x"5653504D", x"4A46423F",
									 -- x"3F3C3A39", x"3836322F", x"2E2A2A2A", x"27272824", x"25252524", x"24232424", x"1F212221", x"2021211F",
									 -- x"1F1F1E1E", x"1D1C1C1B", x"1B1B1B1A", x"19191A1B", x"18171616", x"16161515", x"13141412", x"12131210",
									 -- x"12100F10", x"0E0C0B0C", x"0E0D0C0B", x"0B0C0D0D", x"0B0C0D0D", x"0C0B0B0C", x"0E0E0E0D", x"0C0B0B0B",
									 -- x"0A0B0B0B", x"0B0B0B0B", x"0A0A0A0A", x"0A0A0A0A", x"09090909", x"0909090A", x"0B0A0A0B", x"0C0B0908",
									 -- x"0A0A0A0A", x"0A0A0A09", x"0A0B0B0A", x"090A0907", x"0A090807", x"07080807", x"07090907", x"07080909",
									 -- x"090B0B0A", x"0A0C0C0A", x"0C0B0A0C", x"0C0C0C0E", x"0E0D0C0C", x"0C0C0D0E", x"0B0C0C0C", x"0C0B0C0C",
									 -- x"0E0E0F0F", x"0F0F0F10", x"0F101111", x"1111100F", x"11111111", x"12121211", x"12111011", x"13131211",
									 -- x"13141514", x"13121213", x"14141414", x"15161616", x"17171818", x"19191919", x"1B1C1C1D", x"1D1C1C1C",
									 -- x"1F222524", x"23232220", x"23262223", x"23242927", x"28292B2B", x"2A292B2C", x"2B2C2B2C", x"30303035",
									 -- x"BDC0C2C1", x"C2C3C3C3", x"C1BCBBBF", x"BEB8B7BA", x"BBBAB9B7", x"B5B1AEAB", x"A8A4A1A1", x"A2A2A2A2",
									 -- x"A2A19EA0", x"A6AAA69E", x"9E9D9FA3", x"A5A29F9C", x"9B9A9895", x"93918B85", x"83807C79", x"75727171",
									 -- x"74787B7A", x"756F6D6C", x"6A67625F", x"5D5D5D5D", x"59585756", x"55545353", x"52525252", x"52514F4D",
									 -- x"4C4C4C4B", x"4A4A4B4C", x"4F4C4B4A", x"4A494B4D", x"4E4C4A4B", x"4E4F4F4E", x"4D4C4A4A", x"4D4F4F4C",
									 -- x"4F4F4F4E", x"4E4E4F51", x"585C5B5A", x"5F616163", x"63676A6A", x"696A6B6B", x"69696664", x"67676669",
									 -- x"686A6C6C", x"6A6A6B6C", x"716E6D70", x"72727374", x"70767373", x"74757974", x"75747678", x"7B7F858A",
									 -- x"8B898588", x"91959699", x"9D9FA0A1", x"A5ADB1B1", x"B4B5B4B4", x"B7B5B3B6", x"B2B4B5B5", x"B6BABFC1",
									 -- x"BEBCBDC1", x"C4C4C7CA", x"CED6DCDF", x"E2E3E8F0", x"F0EDEBEA", x"E9E7E6E6", x"EBEDEEEF", x"F3F7F8F6",
									 -- x"EFEFF0F0", x"F0F1F3F4", x"F2F1F0F0", x"F2F4F4F3", x"F6F2F1F6", x"FBFDFCFA", x"F5F4F4F6", x"F8FAF9F8",
									 -- x"FAFCFEFE", x"FDFCFCFD", x"F8F3EFEB", x"E7E5E1D9", x"D1C9C6C8", x"CBCFD2D0", x"D1CDC9C7", x"C7C6C7C9",
									 -- x"C4C4C3BF", x"BBB5AFAC", x"ABACABA5", x"9E97908B", x"827B756E", x"6765615A", x"57555250", x"4E4B4542",
									 -- x"403C3838", x"3938322D", x"2F2A2828", x"26272722", x"25252524", x"23222121", x"1F21211F", x"1E1F2020",
									 -- x"1F1E1E1D", x"1C1C1C1C", x"1B1B1A19", x"18181819", x"19181716", x"15151413", x"13131311", x"11111110",
									 -- x"11101010", x"0F0D0C0D", x"0D0C0B0A", x"0A0B0C0C", x"0D0E0D0D", x"0B0B0B0C", x"0D0E0E0E", x"0D0C0C0B",
									 -- x"0D0C0B0A", x"0A0A0B0C", x"0A0A0A0B", x"0B0A0A09", x"0A0A0908", x"08090A0A", x"0A0A0A0A", x"0B0A0908",
									 -- x"0A0A0909", x"090A0A0B", x"0B0B0A09", x"0A0B0A07", x"0B090807", x"08080908", x"090A0A07", x"07080A09",
									 -- x"090B0B0A", x"0A0B0B0A", x"0C0B0B0C", x"0D0C0C0E", x"0E0E0D0C", x"0C0C0D0D", x"0C0C0C0B", x"0B0B0D0E",
									 -- x"0D0E0F0F", x"0E0E0F10", x"0F101112", x"12111110", x"10100F10", x"11111111", x"11111212", x"13131313",
									 -- x"15151413", x"11111314", x"14141515", x"16171717", x"17181818", x"18191919", x"1C1C1D1D", x"1C1C1C1C",
									 -- x"21232422", x"21222222", x"23262324", x"24242825", x"27282A2A", x"2A2A2B2C", x"2C2C2A2B", x"30302F32",
									 -- x"C1C2C2C0", x"C0C2C4C3", x"C3BFBFC3", x"C3BEBEC4", x"C3C2C1C2", x"C3C4C2C0", x"BAB4AEAC", x"ADADADAD",
									 -- x"B1ACA8A9", x"B0B5B3AC", x"AAA8A9AE", x"B0AFABA8", x"A7A49D96", x"9392908D", x"908D8883", x"7F7B797A",
									 -- x"797C807F", x"7B777676", x"706F6C69", x"66656565", x"65646363", x"62605F5D", x"5B5B5B5C", x"5B595653",
									 -- x"53514E4C", x"4B4C4E4E", x"4D4B4948", x"48474748", x"494A4A48", x"47474A4C", x"4A484747", x"494B4A47",
									 -- x"4C4C4C4C", x"4C4D4E50", x"54585756", x"5B5D5E60", x"5E616261", x"61636565", x"66655E5A", x"5C5E6064",
									 -- x"60626262", x"61606163", x"68656469", x"6F72716F", x"696E6D70", x"71717673", x"72727479", x"7C7E8184",
									 -- x"82858486", x"8B929DAA", x"ABAEAEAA", x"ABB2B6B5", x"B5B4B1B3", x"B6B3B1B5", x"B1B2B3B4", x"B5B8BBBD",
									 -- x"BDBCBDC0", x"C3C5C8CC", x"D1DBE3E9", x"ECEAEBF1", x"F0ECEAEA", x"EAE8E6E6", x"EAECEDEE", x"F2F6F7F7",
									 -- x"F3F1EFEF", x"F0F1F2F3", x"F3F1F0F1", x"F3F4F3F1", x"F5F4F5F9", x"FCFCF9F6", x"EDEEF1F3", x"F4F5F5F5",
									 -- x"F7F7F9FA", x"FAF7F2EF", x"ECE6E0DC", x"D9DBDBD5", x"D2C9C5C5", x"C6C9CCCB", x"C9C6C2C0", x"BEBDBFC1",
									 -- x"C3C1BDB8", x"B3AEAAA8", x"A4A6A49F", x"99948F8B", x"827B746F", x"6966645E", x"5A575452", x"514D4844",
									 -- x"413D3A39", x"3938322D", x"2F2A2828", x"25262723", x"25242322", x"2120201F", x"1E202120", x"1E1E1F20",
									 -- x"201F1D1C", x"1B1B1A1A", x"1A1A1918", x"16161616", x"17161615", x"15151413", x"11121211", x"11111111",
									 -- x"100F0F10", x"100F0E0F", x"0C0C0B0B", x"0B0B0C0C", x"10100F0E", x"0D0D0D0E", x"0C0D0E0D", x"0D0C0C0C",
									 -- x"0E0D0C0B", x"0A0A0B0B", x"0A0A0B0B", x"0B0A0909", x"09090808", x"08090A0B", x"0A0A0A0A", x"0A090808",
									 -- x"09090909", x"090A0A0A", x"0B0B0A09", x"090B0A08", x"0B0A0808", x"08090909", x"0A0A0A08", x"07090A0A",
									 -- x"0A0B0B0A", x"0A0B0B09", x"0A090A0B", x"0C0B0B0C", x"0D0D0C0C", x"0C0C0C0C", x"0C0D0D0C", x"0C0C0D0E",
									 -- x"0D0E0F0F", x"0D0D0E0F", x"0E0F1012", x"12111010", x"100F0E0F", x"10111111", x"10111314", x"13141516",
									 -- x"17161513", x"11111315", x"14141516", x"16171819", x"18181818", x"19191A1A", x"1B1C1D1E", x"1D1D1E1F",
									 -- x"1E202121", x"21222324", x"23262325", x"25242725", x"25272829", x"292A2B2C", x"2D2D2A2B", x"31323031",
									 -- x"C3C4C4C2", x"C2C4C6C6", x"C4C4C4C5", x"C5C5C7C9", x"CBC9C7C7", x"C9CAC9C7", x"C1BBB4B2", x"B3B4B4B5",
									 -- x"BAB7B4B6", x"BBBFBFBC", x"BAB8B7BA", x"BCBBB8B6", x"B3B1AAA1", x"9B9A9B9C", x"9C97928F", x"8B888789",
									 -- x"86868786", x"84828181", x"7C7D7C79", x"76747373", x"73727272", x"716E6A68", x"64646668", x"6A696562",
									 -- x"5C595653", x"5251504F", x"4E4C4A4A", x"4A484748", x"46464644", x"43434548", x"47454546", x"48494847",
									 -- x"4A4A4A4A", x"4A4B4D4E", x"50545353", x"575A5A5C", x"5D5E5D5A", x"585A5C5C", x"5D5F5D5C", x"5D5A5759",
									 -- x"5A5B5B5B", x"5B5B5D5E", x"615F5F64", x"6C706E69", x"6364646C", x"6F6C7275", x"72727377", x"7A7B7D7F",
									 -- x"7B82878A", x"8D919BA8", x"ADB5B9B7", x"B7BABBB8", x"B8B6B3B5", x"B9B6B3B7", x"B3B3B3B5", x"B6B8BBBD",
									 -- x"BDBCBDBF", x"C1C3C8CC", x"D2DCE7F1", x"F6F3EFF1", x"EFECE9E9", x"EAE9E8E9", x"ECEFF0F0", x"F1F3F4F4",
									 -- x"F8F4F0EF", x"F1F3F4F3", x"F4F2F1F2", x"F3F4F3F1", x"EFF1F1F1", x"F1F0EFEE", x"E6EAEEF0", x"EFEEEFF1",
									 -- x"F4F3F2F3", x"F5F2ECE7", x"E3DCD6D3", x"D3D7D8D2", x"CEC7C4C3", x"C0C1C4C4", x"C4C0BDBB", x"B9B7B7B9",
									 -- x"BEBCB9B4", x"AFABA7A5", x"A1A19E99", x"94908D8A", x"837B7570", x"6A676560", x"5D595452", x"514E4A46",
									 -- x"44413F3C", x"3B383432", x"2F2C2B2A", x"25252725", x"24232120", x"20201F1E", x"1B1C1D1E", x"1C1B1B1C",
									 -- x"1D1C1B1A", x"19181818", x"18181817", x"16151516", x"13131314", x"15161615", x"12121313", x"12111112",
									 -- x"100F1011", x"110F0F0F", x"0F0F0E0E", x"0E0E0F0F", x"11110F0F", x"0E0F1010", x"0E0E0E0D", x"0C0C0D0D",
									 -- x"0D0D0C0C", x"0B0A0A09", x"0A0A0B0B", x"0B0B0A09", x"08090909", x"090A0909", x"09090A09", x"09080808",
									 -- x"08080909", x"09090909", x"0A0B0C0A", x"08090A0A", x"0B0A0908", x"09090A09", x"0A0B0A08", x"080A0B0A",
									 -- x"0A0C0C0A", x"0A0B0B09", x"0908090C", x"0C0B0A0B", x"0B0C0C0D", x"0D0D0D0D", x"0B0B0C0C", x"0C0C0D0D",
									 -- x"0E0F100F", x"0E0D0E0E", x"0E0F1011", x"1110100F", x"100F0E0E", x"0F101111", x"11121414", x"14141517",
									 -- x"17171715", x"13131415", x"14151616", x"16171819", x"18181819", x"1A1B1C1C", x"1C1D1F1F", x"1E1E1F20",
									 -- x"1D1F2223", x"23232324", x"23262326", x"27242826", x"28292A2B", x"2C2D2D2E", x"2E2F2D2D", x"32333031",
									 -- x"BFC1C2C1", x"C2C5C6C6", x"C5C7C7C6", x"C7CBCCCB", x"CFCCC9C8", x"C8C9C8C6", x"C1BCB7B7", x"B9BABBBD",
									 -- x"BEBFBFC1", x"C4C6C5C4", x"C4C1BFC0", x"C1BFBEBD", x"BCBDBBB4", x"AEADAEAE", x"ABA6A2A0", x"9C989698",
									 -- x"99989693", x"918F8D8B", x"8C8C8B89", x"86838181", x"807F7E7E", x"7C797471", x"71727376", x"78777470",
									 -- x"69686663", x"5F5B5755", x"53504D4C", x"4B494747", x"48444040", x"43444341", x"41414346", x"47464748",
									 -- x"4B4B4A49", x"494A4B4C", x"4F535352", x"55565556", x"5A5A5956", x"55565858", x"575B5A59", x"59555152",
									 -- x"54555657", x"595A5C5D", x"5D5C5C60", x"686D6A63", x"5F5D5D67", x"69656C72", x"73717173", x"75777B7E",
									 -- x"7E828487", x"8C8E949C", x"A4AFBABF", x"C0C1C1BF", x"BDBCB8B9", x"BDBAB6B6", x"B6B3B2B2", x"B4B7BABE",
									 -- x"BFBFBFBF", x"C0C3C7CB", x"CDD5E1F0", x"FAF9F5F7", x"F3F0EDEB", x"EAEAEDF1", x"EDEFF1F0", x"F1F3F5F6",
									 -- x"F8F6F3F3", x"F4F5F6F5", x"F5F3F2F1", x"F1F0EFED", x"EBECEBE7", x"E4E5E8EB", x"E4E8ECEC", x"EAE9EBED",
									 -- x"F1EEEBEC", x"EEEEEBE7", x"DFD9D4D2", x"D1D5D4CE", x"C8C4C2C1", x"BBBABDBE", x"C2BEBAB8", x"B5B2B1B1",
									 -- x"B8B8B8B6", x"B2ADA8A5", x"A19F9A94", x"908E8B88", x"837A7571", x"6B676460", x"5E5A5451", x"514F4B47",
									 -- x"4544423E", x"3A373635", x"32302F2D", x"27252625", x"24222121", x"2121201E", x"1B1B1B1D", x"1D1B1A1A",
									 -- x"1A1A1A19", x"19191919", x"15161717", x"16161616", x"14141414", x"15141312", x"14141414", x"12101012",
									 -- x"12111112", x"120F0E0E", x"100F0F0F", x"0F101010", x"11100F0E", x"0F101010", x"10100F0E", x"0D0D0E0F",
									 -- x"0D0D0D0C", x"0C0B0A09", x"0A0A0B0B", x"0B0A0A0A", x"0A0A0A0A", x"09090807", x"090A0A09", x"08080809",
									 -- x"08080909", x"09090908", x"080B0C0A", x"0808090A", x"0A090909", x"090A0909", x"090A0A09", x"0A0C0C0A",
									 -- x"0B0C0C0B", x"0B0B0B09", x"09090B0D", x"0E0C0B0C", x"0C0C0D0E", x"0F0F0F0E", x"0C0C0D0E", x"0D0D0E0E",
									 -- x"10101010", x"100F0F0F", x"0F0F0F10", x"100F0F0F", x"0F0F0F0F", x"10111111", x"13141514", x"13121315",
									 -- x"16171717", x"15141415", x"14161717", x"16171819", x"19191919", x"1A1C1D1E", x"1E202222", x"201E1E1F",
									 -- x"1F212527", x"27242324", x"24262327", x"28252928", x"292A2B2C", x"2D2E2F2F", x"3032302E", x"32323030",
									 -- x"BBBDBFBF", x"C0C2C4C5", x"C7C9C9CA", x"CCCFCECC", x"CECCCAC8", x"C7C7C5C4", x"BEBCBABC", x"BEC0C2C5",
									 -- x"C3C4C5C6", x"C6C6C6C6", x"C6C3C2C2", x"C2C1C1C2", x"C3C5C5C2", x"BFBEBDBC", x"BEBBB9B9", x"B6AFADAE",
									 -- x"ACACABA9", x"A5A29E9B", x"9B9A9795", x"928F8D8C", x"8E8D8B8A", x"8A888481", x"83838487", x"89888581",
									 -- x"7F7D7B77", x"726D6A68", x"635D5753", x"504C4949", x"4B474241", x"4343413D", x"3D3E4144", x"43414245",
									 -- x"47484849", x"4849494A", x"4E52514F", x"52525050", x"53545453", x"53555655", x"56575450", x"504E4E51",
									 -- x"4E4F5153", x"5558595B", x"5859585A", x"6269665E", x"5D5D5A60", x"605D6468", x"6D6C6D70", x"7274787C",
									 -- x"80817F80", x"85888C93", x"98A2AFB7", x"BBBEC3C6", x"C8C8C4C3", x"C6C5BFBC", x"BAB7B4B4", x"B5B7BABE",
									 -- x"C1C2C2C2", x"C2C4C8CB", x"CED4DDEA", x"F5F6F5F9", x"F7F4F0EB", x"E6E7EDF5", x"F0F1EFEE", x"F0F3F4F4",
									 -- x"F1F3F5F6", x"F5F5F6F7", x"F7F5F2EE", x"EAE6E4E2", x"E7E9E7E2", x"DFE3E9ED", x"E2E3E3E3", x"E2E3E4E5",
									 -- x"E9E7E5E5", x"E6E6E4E3", x"DDD9D6D3", x"D0D1D0CB", x"C5C1C0BF", x"B9B8BABB", x"BEBBB9B7", x"B2AEADAE",
									 -- x"B1B2B1B0", x"ACA8A3A1", x"9D99938D", x"8B8A8783", x"81787370", x"6B676460", x"5E595451", x"51504C49",
									 -- x"4847433F", x"3B383737", x"3632312F", x"2A282825", x"24232323", x"2423201D", x"1F1C1B1D", x"1E1D1C1C",
									 -- x"1A1A1A1B", x"1A1A1A1A", x"14151718", x"17151414", x"16161515", x"1412100F", x"14131414", x"120F0F12",
									 -- x"12121213", x"120F0E0E", x"0F0F0F0F", x"0F0F0F10", x"11100F0F", x"10101010", x"1011100F", x"0E0D0E0E",
									 -- x"0D0D0D0D", x"0C0B0B0A", x"0B0B0B0B", x"0B0A0A0A", x"0B0A0A09", x"09080808", x"090A0A09", x"08080809",
									 -- x"09090808", x"08080808", x"080A0A09", x"09090908", x"09090909", x"0A0A0908", x"08090A0A", x"0B0D0D0B",
									 -- x"0C0D0D0C", x"0B0C0B0A", x"0A0A0C0E", x"0F0D0C0C", x"0C0D0E0F", x"0F0F0E0E", x"0E0E0E0E", x"0E0E0F11",
									 -- x"100F0E0F", x"1111110F", x"1010100F", x"0F0F0F0F", x"100F1010", x"12121211", x"14141312", x"11111213",
									 -- x"15161717", x"15141415", x"15171818", x"1717181A", x"1A1A1A1A", x"1B1D1E1F", x"1E212424", x"211F1F20",
									 -- x"21222629", x"28242223", x"25262328", x"29262A2A", x"292A2A2C", x"2D2E2E2E", x"2F33312F", x"32323031",
									 -- x"BEC0C0C0", x"C1C3C5C5", x"CBCBCCCF", x"D3D3D1CF", x"CFCECCC9", x"C6C4C1C0", x"BCBBBCBE", x"C0C2C4C7",
									 -- x"C8C7C5C4", x"C4C5C6C7", x"C5C4C3C5", x"C5C5C6C8", x"C7C7C7C5", x"C4C5C4C2", x"C1BFC0C4", x"C3BDBBBC",
									 -- x"B9BBBCBB", x"B8B3AFAC", x"B2AFABA7", x"A4A2A09E", x"9B999797", x"97979593", x"90909196", x"999A9895",
									 -- x"928F8B85", x"807D7D7E", x"756D645C", x"57514E4D", x"4E4D4A46", x"42403F3E", x"3B3D4042", x"3F3C3D41",
									 -- x"40424445", x"46464647", x"4A4E4C4A", x"4D4D4A4B", x"4E505150", x"4F4F4E4C", x"5153504D", x"4D4B4A4D",
									 -- x"4B4C4E50", x"52545556", x"54545455", x"5D65645D", x"5D5F5B5A", x"59575E5F", x"6264686C", x"6F707377",
									 -- x"797E8082", x"8584878E", x"9399A2AB", x"B0B6C0CA", x"D5D7D3D1", x"D4D4CDC7", x"C1BDBBBB", x"BBBBBCBE",
									 -- x"C0C2C4C4", x"C4C7CACD", x"D9DCE0E7", x"EEEDEDF4", x"F5F3EEE6", x"E0E0E9F3", x"F9F5F0EC", x"EDEFEEEC",
									 -- x"E8EEF5F7", x"F5F3F5F7", x"F9F6F1EA", x"E3DCD9D7", x"D9DBDAD7", x"D6DAE0E2", x"DEDBD8D7", x"D8DADBDB",
									 -- x"DFE0E1E1", x"DFDDDBDB", x"DBD9D7D4", x"CECDCDC9", x"C3BEBDBD", x"B8B7B9B9", x"B8B8B7B5", x"B0ABABAD",
									 -- x"AAA9A6A3", x"9F9C9998", x"96928B86", x"8585827E", x"7E757170", x"6B676461", x"5D595452", x"52514D49",
									 -- x"4D4A4641", x"3E3C3B3B", x"37323130", x"2D2C2B26", x"24242526", x"2725201D", x"211C191B", x"1D1D1C1C",
									 -- x"1A1A1A1A", x"19181717", x"15171819", x"17141211", x"12121314", x"14141312", x"12121314", x"120F1013",
									 -- x"11111213", x"13100F0F", x"10101011", x"11111111", x"12111010", x"11111110", x"0F101010", x"0E0D0C0C",
									 -- x"0E0E0E0D", x"0C0C0C0C", x"0B0B0B0A", x"0A0A0A0B", x"0A0A0908", x"0809090A", x"0A0A0A0A", x"0808090A",
									 -- x"0A090807", x"07070809", x"08090908", x"0A0B0906", x"0808090A", x"0A0A0908", x"08090A0A", x"0C0E0D0B",
									 -- x"0D0E0E0C", x"0C0C0C0A", x"0A0A0C0F", x"0F0D0C0C", x"0B0C0D0E", x"0E0E0D0C", x"0D0D0C0B", x"0B0C0E10",
									 -- x"0F0D0C0D", x"1012110F", x"12111010", x"0F0F0F0F", x"10101011", x"12131212", x"13121110", x"10111213",
									 -- x"14151616", x"15141415", x"16181A19", x"1817191A", x"1C1B1B1B", x"1B1D1E1F", x"1D202425", x"23212121",
									 -- x"20222529", x"28242223", x"26272428", x"29262A2A", x"2A2A2B2C", x"2E2E2F2E", x"2D32312F", x"31323132",
									 -- x"C1BFBEC1", x"C4C6C5C4", x"CACCCED0", x"D0CFCECD", x"D2CCC9CA", x"C9C5C2C2", x"BDBCBCBD", x"BFC3C6C9",
									 -- x"C9C9CACA", x"C8C4C4C7", x"C2C3C4C5", x"C5C5C6C7", x"C4C7C8C5", x"C3C4C6C6", x"C4C4C2C1", x"C2C3C2C0",
									 -- x"BFBFBEBE", x"BEBDBBB9", x"BCBAB7B5", x"B4B3B2B2", x"ADAAA6A5", x"A7A9AAA9", x"A7A8A9A8", x"A8A7A8A9",
									 -- x"A19D9A97", x"918A8889", x"857F776E", x"66605B58", x"5154534C", x"46454442", x"403F3E3E", x"3D3D3D3E",
									 -- x"3F3F4041", x"43444546", x"48464347", x"4D4C494D", x"49484A4D", x"4C49494C", x"4C4E4E4D", x"4C4E4D4B",
									 -- x"4D4D4D4D", x"4F515354", x"524F4D4F", x"565C5F60", x"6161605B", x"5655585D", x"5B616061", x"67696E7B",
									 -- x"7F7B8084", x"80848D91", x"93949AA2", x"AAB4C0CA", x"DEE4E7DF", x"D7D8D5CA", x"C4C1C0C0", x"BFBDBEC1",
									 -- x"C2C3C4C7", x"CACED0D0", x"DEE0DEEA", x"F3ECE5DF", x"E0E0E2E2", x"E2EAF4F6", x"F6F7F2EB", x"EBEEE8DD",
									 -- x"D8E6F1F0", x"E8E6EBF1", x"F2F4F0E5", x"DCDADAD8", x"D6D0CED1", x"D4D4D7DD", x"DDDBD7D3", x"D0D0D2D5",
									 -- x"D4D7DAD9", x"D8D8D8D7", x"D5D5D3CF", x"CAC6C4C4", x"BFBCBAB9", x"B7B4B2B2", x"B1B2B4B5", x"B5B2ADAA",
									 -- x"A7A6A29D", x"9B98938D", x"8B888583", x"7F7A7777", x"76706E6B", x"6665635E", x"58575655", x"53504B48",
									 -- x"4D4B4744", x"413F3D3B", x"38393631", x"2F2F2D29", x"27292825", x"2425221E", x"211E1C1C", x"1E1E1D1B",
									 -- x"1A19191A", x"1B191717", x"19171514", x"14151719", x"12121214", x"15151412", x"14131314", x"13111114",
									 -- x"10121213", x"14100D10", x"0E101111", x"1313100D", x"12111111", x"13131211", x"12121210", x"0F0E0F10",
									 -- x"100F0E0F", x"0E0C0A0A", x"0D0C0B0A", x"0A0A0B0B", x"090B0A08", x"07090908", x"0A090909", x"0A090706",
									 -- x"09090909", x"08080809", x"0A0A0909", x"09090909", x"090A0B0A", x"09090A0B", x"090A0A0A", x"0B0D0D0C",
									 -- x"0E0E0D0C", x"0A0A0A0A", x"0D0D0D0D", x"0D0D0D0D", x"0E0E0E0E", x"0D0C0B0A", x"0D0D0D0D", x"0C0D0F11",
									 -- x"0F0D0D10", x"11100F0F", x"110E0D0F", x"10100F0F", x"10111213", x"1312110F", x"10101111", x"12121111",
									 -- x"13121316", x"16141517", x"16171717", x"181A1A18", x"1B1C1A19", x"1D1E1C1D", x"1E222423", x"2221201E",
									 -- x"22232221", x"22242524", x"23262A2B", x"2928292A", x"2B2A2A2C", x"2B2C2F34", x"312F3033", x"33303134",
									 -- x"C5C4C5C7", x"CACBC9C8", x"C9CACCCE", x"CFD0CFCF", x"CECAC8C7", x"C6C5C3C3", x"C1C1C1C2", x"C4C7C8C9",
									 -- x"C9C8C9C9", x"C7C5C5C7", x"C2C3C5C6", x"C6C6C6C6", x"C4C7C7C4", x"C3C4C5C4", x"C4C4C3C2", x"C3C4C3C1",
									 -- x"C1C0C0BF", x"BFBEBCBB", x"BDBCBABA", x"B9B8B6B5", x"B1B0AEAF", x"B0B0AEAB", x"ADAEAFAE", x"ABA9AAAB",
									 -- x"A79F9591", x"8F8D8A87", x"85817B75", x"706C6865", x"5F5D5954", x"514F4C4A", x"46444140", x"40403E3D",
									 -- x"3C3D3D3F", x"41434546", x"484A4745", x"49494747", x"4647494A", x"48464749", x"4C4E4F4F", x"4F4F4E4C",
									 -- x"4D4E5051", x"52515151", x"4F4E4D4F", x"53585C5E", x"5E5E5D5B", x"59575656", x"585D5D5E", x"63656B77",
									 -- x"7A7B8185", x"84868D91", x"979498A2", x"A8ADB8C5", x"CEDDE7E2", x"DDDFDCD0", x"C9C9C7C4", x"C2C3C4C4",
									 -- x"CAC5C4CA", x"D2D6D5D3", x"DCE4DFE0", x"E8EEF0EA", x"DBD8D9DD", x"E2ECF2F0", x"F0EEEBE8", x"E5E1DBD7",
									 -- x"D5DEE4E1", x"DBDBE1E6", x"EBEFEBE1", x"DCDFDDD6", x"D3D0CED0", x"D1D2D5DA", x"D9D8D5D2", x"CFCDCDCE",
									 -- x"CFD2D4D4", x"D3D3D1D0", x"CFCDCAC7", x"C5C2BFBD", x"BBB8B5B4", x"B2AFAFB0", x"AEAEAFAF", x"AFACA7A3",
									 -- x"9F9E9B97", x"95928C86", x"8783807E", x"7C777575", x"746E6C6A", x"6563615D", x"5A585452", x"51504E4D",
									 -- x"4B484543", x"42413E3C", x"39383633", x"31302F2D", x"292A2A28", x"28282624", x"22222121", x"201F1E1D",
									 -- x"1B1A1A1C", x"1C1A1818", x"1A1A1A1A", x"19181717", x"18171616", x"17161412", x"16151516", x"15121112",
									 -- x"14141113", x"16131012", x"10111313", x"1414120E", x"10100F10", x"12131312", x"11111010", x"10101010",
									 -- x"13100E0D", x"0D0C0C0D", x"0D0D0C0C", x"0B0B0A0A", x"0A0B0A09", x"080A0A08", x"0A0A0909", x"0A090806",
									 -- x"09090909", x"08070809", x"09090909", x"0A0A0B0B", x"090A0A09", x"0808090A", x"0A0B0B0A", x"0B0D0E0D",
									 -- x"0F0F0E0D", x"0C0C0C0D", x"0D0E0E0E", x"0E0E0D0D", x"0E0F0F0F", x"0F0E0D0D", x"0E0E0F0F", x"0F101011",
									 -- x"0F0E0E10", x"11100F0E", x"0E0E0E10", x"100F1012", x"10101113", x"13131110", x"11111112", x"12121213",
									 -- x"13131417", x"18161617", x"16191B1B", x"1B1C1C1A", x"1B1C1B1B", x"1F1F1E21", x"1F222322", x"21232322",
									 -- x"23242423", x"24262828", x"25272829", x"29292A2B", x"2D2C2C2D", x"2C2C2E32", x"2E2F3132", x"32343535",
									 -- x"C9CACCCE", x"CFCFCECD", x"CFCFCFCF", x"CFCFCFCF", x"CFCECCC8", x"C7C8C8C8", x"C8C8CACB", x"CDCECDCC",
									 -- x"CAC9C8C8", x"C7C6C5C6", x"C2C3C4C5", x"C5C5C4C5", x"C5C6C5C3", x"C3C3C3C2", x"C3C4C4C3", x"C3C4C3C1",
									 -- x"C2C1C1C0", x"C0BFBEBC", x"BABABBBB", x"BBB9B7B5", x"B3B1B0B1", x"B2B2AFAD", x"AFB0B1AF", x"ABA9A8A9",
									 -- x"A79F958F", x"8F8F8B87", x"8885817E", x"7A777370", x"6D665F5D", x"5C595551", x"4D494442", x"4343413E",
									 -- x"3E3E3F40", x"42444647", x"484D4A45", x"46484644", x"46494B49", x"4747484A", x"4C4E5051", x"52535250",
									 -- x"51525354", x"54545352", x"51515252", x"5355595C", x"59585758", x"58585553", x"54595A5B", x"5E606772",
									 -- x"7A808487", x"89898D94", x"9B9AA1AF", x"B4B1B4BD", x"C8CBCDD6", x"EAF6E8CE", x"CBCBC9C5", x"C4C5C8C9",
									 -- x"CACBD1D6", x"D5D2D5DC", x"DEE7E2E1", x"E6EAEEEA", x"DED8D7DB", x"E2EAEBE5", x"E6E1E2E5", x"E3DBD8DA",
									 -- x"DBE2EAEB", x"E8E4E2E1", x"DFE6E4DD", x"DFE6E3D8", x"D3D3D2D1", x"D1D1D3D5", x"D3D4D4D2", x"D1CECCCA",
									 -- x"CCCECFCE", x"CFCFCCC9", x"C8C4C0BE", x"BFBDB8B4", x"B7B3B0AD", x"AAA8A8AA", x"A7A6A5A6", x"A6A49F9B",
									 -- x"9A989490", x"8E8B8782", x"817D7978", x"76747270", x"706B6967", x"6361605B", x"5B585452", x"51504F4D",
									 -- x"4B494644", x"4442403E", x"3C393635", x"34313031", x"2D2B2B2C", x"2C2A2828", x"21222323", x"211F1E1E",
									 -- x"1D1C1D1E", x"1E1B1918", x"1B1B1C1C", x"1B1A1918", x"17161516", x"17171514", x"16161717", x"16131212",
									 -- x"15141010", x"15131011", x"0F111212", x"1313110E", x"12111011", x"11121212", x"100F0E0F", x"10111110",
									 -- x"13100D0C", x"0C0C0C0E", x"0D0D0D0D", x"0C0B0A09", x"0A0B0B0A", x"090A0A09", x"0B0B0A0A", x"0A090807",
									 -- x"09090909", x"08070809", x"0A0A0A0A", x"0A0B0B0B", x"0A0A0A0A", x"09090A0A", x"0B0C0C0B", x"0C0E0F0E",
									 -- x"0E0E0E0D", x"0D0D0E0F", x"0E0F1010", x"100F0E0D", x"0F0F0F10", x"10101010", x"11100F10", x"11111212",
									 -- x"100F0F11", x"12100E0E", x"0E0F1011", x"100F1114", x"10111213", x"14141311", x"13121212", x"12131414",
									 -- x"14141519", x"1B1A1716", x"171B1F1F", x"1F1F1E1C", x"1A1D1B1B", x"1D1E1E21", x"24252422", x"21212221",
									 -- x"23252624", x"2427292A", x"28272727", x"292A2B2B", x"2C2C2D2E", x"2D2C2E31", x"2F343431", x"30333431",
									 -- x"CBCDD0D1", x"D1D0D0D1", x"D3D3D2D2", x"D1D0CFCE", x"D2D4D1CB", x"C8CACBCA", x"CBCBCCCE", x"D0D1D0CE",
									 -- x"CCCAC8C7", x"C7C6C5C5", x"C1C2C2C2", x"C2C1C2C2", x"C4C4C3C2", x"C3C3C3C2", x"C1C3C3C3", x"C3C3C2C0",
									 -- x"C1C1C0BF", x"BFBEBDBC", x"B8B9B9BA", x"BAB8B6B4", x"B3B0ADAC", x"AEAFAFAF", x"AFAEACAA", x"A9A8A7A7",
									 -- x"A1A09C96", x"92908D8A", x"89878482", x"807E7B78", x"776E6767", x"67635D59", x"55524D49", x"49494643",
									 -- x"45454647", x"48494949", x"4A4E4C48", x"48484748", x"484D4F4C", x"4A4C4E4F", x"50525456", x"58595959",
									 -- x"57575756", x"57575859", x"58585857", x"5757585A", x"59575656", x"595A5958", x"575A5C5D", x"5E606871",
									 -- x"7F878888", x"8C8C8F99", x"9899A1AC", x"B0ACABAD", x"B0B5BAC2", x"D0D8D1C7", x"C8C6C4C4", x"C4C6CCD3",
									 -- x"D4D3D5D4", x"CBC5CFDE", x"E1E3DEE2", x"E4E0E2E4", x"E3DCDADC", x"DFE4E3DE", x"DDD9DADF", x"DFDAD8DB",
									 -- x"D8E0EAF1", x"F2EEE6E0", x"DCE1E1DE", x"E0E5E2D9", x"D7D7D5D2", x"D2D2D1CE", x"CCCDCFD0", x"D0D0CCC9",
									 -- x"C8C9CACA", x"CBCCC9C6", x"C1BEBBBB", x"BBB8B2AD", x"B0ACA8A4", x"A19D9D9E", x"9E9C9B9C", x"9E9D9995",
									 -- x"97938D89", x"87858381", x"7E797472", x"72716E6C", x"6B676665", x"61605F5A", x"5A585654", x"52504D4A",
									 -- x"4A494745", x"43413E3D", x"3F3A3737", x"36323132", x"2F2C2B2D", x"2D292728", x"21212222", x"22212020",
									 -- x"1F1E1E20", x"1F1C1A19", x"1C1B1A19", x"191A1B1C", x"17161516", x"17171615", x"16161717", x"16141414",
									 -- x"14151211", x"14131011", x"10111212", x"1213120F", x"14141312", x"12111111", x"100F0D0E", x"1011100F",
									 -- x"100E0D0E", x"0E0C0B0C", x"0D0D0D0D", x"0C0B0A0A", x"0B0B0B0B", x"0B0B0A0A", x"0C0C0C0C", x"0B0A0808",
									 -- x"090A0909", x"08080809", x"0C0B0B0A", x"0A0A0A0A", x"0B0B0B0A", x"0A0A0B0B", x"0B0C0C0B", x"0B0D0F0F",
									 -- x"0D0E0E0D", x"0D0D0E0F", x"0F101011", x"1110100F", x"0F101011", x"11121212", x"14110F0E", x"10121313",
									 -- x"12100F11", x"12111010", x"11101112", x"11101113", x"12121314", x"15151312", x"13131212", x"12131415",
									 -- x"16151619", x"1B1C1917", x"181D2020", x"1F1F1F1E", x"1D201F1D", x"1E1D1C20", x"26252422", x"21212121",
									 -- x"22252624", x"24262829", x"27282828", x"292A2B2C", x"2A2B2D2E", x"2E2F3032", x"31343431", x"3031312F",
									 -- x"CCCED0D1", x"D0D0D1D3", x"CFD0D1D2", x"D2D1D1D0", x"D1D2CFCA", x"C7C9CAC8", x"C8C7C8CA", x"CCCDCDCC",
									 -- x"CCCBC9C7", x"C6C5C4C3", x"C2C2C1C0", x"BFBFC0C1", x"C2C1C0C1", x"C1C1C1C1", x"C1C3C3C2", x"C2C2C2C0",
									 -- x"C0C0BEBE", x"BEBDBCBC", x"BABAB9B9", x"B8B7B6B5", x"B5B1ADAC", x"ADAEAFAF", x"AFABA7A6", x"A8A9A8A7",
									 -- x"A3A3A09C", x"98969390", x"8B898786", x"86858382", x"7E777273", x"736D6764", x"605F5A54", x"504F4E4B",
									 -- x"4A4B4D4E", x"4E4E4D4C", x"4D4F4D4D", x"4D49484E", x"4B505250", x"4F525454", x"5758595B", x"5C5E5F60",
									 -- x"5C5C5B5A", x"5A5B5C5C", x"5D5C5B5A", x"5A5A5A59", x"5C5C5D5E", x"5F606263", x"61616365", x"63656C72",
									 -- x"7F888B8B", x"8F90939C", x"9A9C9E9F", x"A1A4A4A3", x"A4ADB3B7", x"BBB9BBC4", x"C8C3C2C7", x"C8C8D2DF",
									 -- x"E7D6C8C4", x"C6C9D2DD", x"E5E4DCDE", x"E1DDE0E3", x"DFDBDCDC", x"DBDCDFDE", x"DBD8D5D5", x"D6D5D3D2",
									 -- x"D5D9DFE6", x"EBEBE8E6", x"DEDFDFDE", x"DDDAD7D5", x"D5D3D1CF", x"CFCFCBC5", x"C4C6C9CB", x"CECFCCC8",
									 -- x"C5C6C6C6", x"C7C8C6C2", x"BDBCBBBA", x"B8B4AEA9", x"A5A29E9B", x"97939192", x"96949394", x"96959390",
									 -- x"908C8784", x"82807D7C", x"7B777370", x"6F6E6C69", x"67646565", x"615F5E5B", x"5A585554", x"52504D4A",
									 -- x"46474846", x"423E3D3D", x"413D3939", x"37323032", x"302D2C2E", x"2D292728", x"26242222", x"23242221",
									 -- x"201F1F20", x"201D1A1A", x"1D1C1A18", x"181A1C1D", x"1C1A1918", x"18171614", x"16171715", x"14151516",
									 -- x"15181715", x"15131113", x"12141514", x"14141412", x"14141413", x"12111111", x"110F0E0F", x"1111100E",
									 -- x"100E0E0F", x"0F0E0D0D", x"0E0D0D0C", x"0C0C0C0D", x"0C0B0C0C", x"0C0B0B0B", x"0D0D0D0D", x"0C0A0A09",
									 -- x"0A0A0A09", x"09080909", x"0C0B0B0A", x"0A090909", x"0B0B0A0A", x"0A0B0B0B", x"0B0D0D0B", x"0B0D0E0F",
									 -- x"0F0F0F0E", x"0D0D0E0F", x"10101010", x"10111213", x"10101111", x"12121213", x"14121111", x"12131312",
									 -- x"14110F10", x"12121213", x"13101011", x"12121112", x"14141415", x"15151413", x"13131212", x"13141515",
									 -- x"17161617", x"1A1C1B19", x"1A1E201F", x"1E1F2020", x"21242321", x"22201F22", x"21212122", x"23232425",
									 -- x"23262625", x"24262727", x"25282A2A", x"29292B2D", x"2B2D2E2F", x"30323333", x"2F2E2F32", x"32303033",
									 -- x"CECFD0D0", x"D0D0D1D2", x"D0D1D1D2", x"D2D1D0D0", x"CDCDCCC9", x"C8C9C9C9", x"C8C6C4C5", x"C8CACAC9",
									 -- x"C9C9C8C5", x"C4C3C2C1", x"C2C2C1C0", x"BFBEBFC0", x"BEBDBDBE", x"BFBEBEC0", x"C0C2C2C1", x"C0C0C0BF",
									 -- x"BFBDBCBC", x"BBBBBBBA", x"BAB8B6B5", x"B4B4B3B3", x"B2B0AEAD", x"AEADACAA", x"ACA8A4A3", x"A5A7A6A5",
									 -- x"A9A29C9B", x"9B999694", x"94928F8E", x"8C8B8886", x"817E7B7B", x"7B77716D", x"6968635B", x"5554524F",
									 -- x"4E4F5153", x"54535251", x"54535151", x"514C4A50", x"4E515353", x"54565758", x"5B5A5A5C", x"5D5D5E60",
									 -- x"5E5F5F60", x"5F5F5E5E", x"605E5D5E", x"5F5F5F5E", x"6164686A", x"6B6C6E70", x"706C6D6E", x"6A6C7173",
									 -- x"7B858C8D", x"8F92979D", x"9FA4A6A5", x"A5A8A39C", x"AAACACB6", x"C8CCCBD1", x"D0CBCCD0", x"CFCDD7E4",
									 -- x"E3D4C9CC", x"D5DCE2E6", x"ECF4EEEA", x"EAE9E9E2", x"DFDDDEDD", x"D8D7DCDD", x"DBDAD6D2", x"D3D6D4D1",
									 -- x"D9DBE0E4", x"E5E4E3E4", x"DBD8D7D8", x"D4CFCDD0", x"CCC9C7C7", x"C8C6C2BE", x"C0C3C6C9", x"CED2CFC9",
									 -- x"C7C8C7C5", x"C4C3C2BF", x"BABABAB8", x"B4AEA9A5", x"9E9B9997", x"948F8D8D", x"8E8E8D8D", x"8D8C8A88",
									 -- x"88858382", x"807C7875", x"7775716E", x"6D6D6A67", x"66646565", x"615F5E5B", x"5A585452", x"51504F4E",
									 -- x"48494A49", x"46434141", x"423F3C3B", x"38353332", x"302E2E2E", x"2E2C2A2A", x"29262322", x"2323211E",
									 -- x"21201F20", x"201D1B1B", x"1D1D1D1C", x"1C1B1B1B", x"19181818", x"18181715", x"18191715", x"14151616",
									 -- x"14191916", x"15131114", x"12141514", x"13141413", x"12131413", x"13121212", x"12111011", x"1212100F",
									 -- x"14110F10", x"10101012", x"0F0E0E0D", x"0D0E0E0F", x"0D0D0D0F", x"0F0D0D0D", x"0D0D0E0E", x"0C0B0B0B",
									 -- x"0B0B0B0A", x"09090A0A", x"0A0A0A0A", x"0A0A0A0B", x"0B0A090A", x"0A0B0A0A", x"0B0D0D0B", x"0A0C0E0F",
									 -- x"11111110", x"0F0F0F10", x"11101010", x"11121415", x"11111111", x"12121313", x"13131516", x"17151311",
									 -- x"15121011", x"12121314", x"120F0E11", x"13131313", x"15151515", x"15151312", x"13131313", x"13141516",
									 -- x"17171616", x"181C1D1C", x"1C1E1F1E", x"1E1F2121", x"21242322", x"24232123", x"21202123", x"24242424",
									 -- x"26272726", x"26272725", x"24282B2C", x"2A292B2E", x"2E303030", x"31323332", x"2F2D2E32", x"322E2F33",
									 -- x"CECFD0D0", x"CFCECECE", x"CFCFCFCE", x"CECDCDCD", x"CCCAC9CA", x"CBCAC9C9", x"CAC7C4C4", x"C6C7C6C5",
									 -- x"C4C6C6C4", x"C1C1C1C0", x"C1C1C1C0", x"BFBDBDBD", x"BBBABBBC", x"BBB9BABD", x"BDBFBFBD", x"BBBBBBBB",
									 -- x"BBB9B8B7", x"B7B7B7B6", x"B5B4B1B0", x"AFAFAFAF", x"ADACABAB", x"ACACA9A6", x"A9A7A5A3", x"A2A1A1A0",
									 -- x"A49B9595", x"94908F91", x"98979593", x"92908C8A", x"84817E7D", x"7F7F7972", x"6F6E6860", x"5B5B5954",
									 -- x"54555758", x"59595959", x"5A5B5856", x"56525053", x"54545558", x"5A5A5B5C", x"5C5B5C5E", x"5F5E5F61",
									 -- x"61616263", x"64646565", x"67686868", x"6868696A", x"6D707578", x"7C7F8387", x"867F7E7E", x"78787C7A",
									 -- x"7E848C8D", x"8C929CA0", x"A1A8AFB3", x"B3AFA398", x"9FACAFB5", x"C6D0D6E2", x"E1E2E1DE", x"D8D7DCE2",
									 -- x"DADCE0E4", x"E6E7EBEF", x"F3FFFCF6", x"F2ECE9E1", x"E1DDDDDC", x"D7D5D8D8", x"D9D9D6D3", x"D3D5D6D5",
									 -- x"D5D9DFE2", x"DFD9D8D9", x"D5D3D0CD", x"CAC7C8CA", x"C3C1C0C2", x"C1BCB9B9", x"BBBFC4C9", x"D0D6D3CD",
									 -- x"CCCCC9C4", x"BFBDBBB9", x"B6B5B3B0", x"ADA8A4A1", x"9B989694", x"918C8A8A", x"87878786", x"85838180",
									 -- x"827E7C7C", x"7A767270", x"71716F6C", x"6B6C6B68", x"67656767", x"625F5E5A", x"5B595554", x"5352504F",
									 -- x"4D4C4C4C", x"4B484542", x"40403E3C", x"3A393734", x"3031302E", x"2E2E2C29", x"27262423", x"22211F1E",
									 -- x"22202020", x"201E1D1D", x"1C1D1E1E", x"1D1C1A19", x"16161617", x"19191817", x"17191816", x"15171817",
									 -- x"13181713", x"14141314", x"12141413", x"12131413", x"13141616", x"15141414", x"13131414", x"13131212",
									 -- x"14121112", x"12121213", x"11101010", x"10101010", x"0F0E0F11", x"110F0F10", x"0C0E0F0E", x"0D0C0C0C",
									 -- x"0B0C0C0B", x"0A0A0A0B", x"0B0B0B0A", x"0A0B0B0B", x"0C0B0A0B", x"0C0C0C0B", x"0C0E0E0C", x"0B0C0F10",
									 -- x"12121110", x"100F1011", x"11111011", x"11121314", x"12121212", x"12131415", x"13151617", x"16151413",
									 -- x"14111011", x"12121112", x"110F0F11", x"12121214", x"14141314", x"14141312", x"13131414", x"15151616",
									 -- x"17181817", x"181C1E1D", x"1D1F1F1F", x"1F212221", x"1F222222", x"25242121", x"25222224", x"25242324",
									 -- x"27272727", x"28292723", x"26282A2B", x"2B2B2C2D", x"2F30302E", x"2F31312F", x"2F2F3031", x"30303031",
									 -- x"CDCECFCF", x"CFCDCBC9", x"C7C7C7C7", x"C8C9CACB", x"CBC7C6CA", x"CCC9C7C7", x"CAC7C4C3", x"C4C4C2C0",
									 -- x"C0C4C5C2", x"C0BFC0BF", x"BEBFC0C0", x"BFBCBBBA", x"B9B9BABA", x"B8B6B7BB", x"B9BBBBB8", x"B6B6B7B6",
									 -- x"B7B6B4B3", x"B3B3B3B3", x"B3B1AFAE", x"AEAEADAD", x"AAA8A8A9", x"ABABAAA8", x"A8A9A8A5", x"A19E9D9E",
									 -- x"98939191", x"8A82848C", x"92929395", x"9695928F", x"8784807F", x"82857F76", x"75726C64", x"6364615C",
									 -- x"5C5C5C5D", x"5D5E5F60", x"5D615E58", x"59595755", x"5A58595D", x"605E5E5F", x"5F5E6063", x"65646566",
									 -- x"64646363", x"65696D6F", x"71737473", x"71707275", x"7C7D8084", x"8A929A9E", x"9B91908F", x"87868984",
									 -- x"85868C8B", x"8791A0A4", x"ADB0B7BE", x"BFB8ACA4", x"A1B2B4B0", x"BCC9D1DC", x"F2F8F7EB", x"E2E1E2E1",
									 -- x"E4EAF0EE", x"E8E5E7EB", x"F5F9F4F2", x"EBE0E1E5", x"DDD7D6D8", x"D6D5D5D3", x"D5D5D3D1", x"CFCED0D2",
									 -- x"D0D5DBDD", x"D9D4D7DC", x"D7D5CFC7", x"C2C2C2C0", x"C0BEBFC2", x"BDB6B4B8", x"B5BAC0C7", x"D0D7D5CF",
									 -- x"CECDC9C1", x"BAB6B3B1", x"B3B1ADA9", x"A7A4A09D", x"99969390", x"8C888585", x"81828382", x"807D7C7C",
									 -- x"7E787372", x"716E6C6C", x"6D6E6E6B", x"6A6B6B69", x"69676968", x"625F5D59", x"5B595857", x"56534F4C",
									 -- x"504D4A4A", x"4B49433E", x"3E403F3C", x"3B3C3A36", x"3233322E", x"2D2D2B27", x"26272827", x"25232121",
									 -- x"23212020", x"201F1E1F", x"1B1B1C1C", x"1C1C1B1B", x"1A19191A", x"1B1A1816", x"15181917", x"17191A19",
									 -- x"16191613", x"16171617", x"14161614", x"13141515", x"16181919", x"18161515", x"14151616", x"15141414",
									 -- x"11101214", x"15131110", x"12121212", x"1211100F", x"11101113", x"13111011", x"0C0E0F0F", x"0E0D0D0D",
									 -- x"0C0C0C0B", x"0B0A0B0B", x"0D0D0C0B", x"0B0A0A0A", x"0F0D0C0D", x"0E0E0E0D", x"0D0F0F0C", x"0B0D1011",
									 -- x"10111010", x"0F0F1011", x"11111112", x"12121313", x"12121212", x"13141516", x"15151513", x"12121416",
									 -- x"13111012", x"13110F0F", x"11111112", x"110F1114", x"13121212", x"13131312", x"14141515", x"16161717",
									 -- x"16191918", x"191C1E1E", x"1E202020", x"21232321", x"21232324", x"28262221", x"24212023", x"25252628",
									 -- x"26262627", x"292A2622", x"2728292A", x"2B2C2D2D", x"2D2E2D2B", x"2C2E2F2D", x"2A2E302F", x"30343533",
									 -- x"CCCECFD0", x"CECBCBCB", x"C8C3C4C6", x"C3C3C7C8", x"C8C9C9C9", x"C9C8C7C7", x"C7C4C2C3", x"C3C0BFC0",
									 -- x"C0C1C1C0", x"BFBFBFBD", x"BFBFBEBE", x"BEBCBAB8", x"BBB7B4B4", x"B5B5B6B7", x"B4B5B6B5", x"B3B2B5B7",
									 -- x"B3B2B3B4", x"B0ABABAF", x"ADADAEAE", x"AEADACAC", x"AAA9A8A8", x"A8A8A9A9", x"AAA7A5A4", x"A5A4A19E",
									 -- x"9C938C89", x"8785878B", x"8C8A8889", x"9096958F", x"8986807E", x"83888680", x"7D787370", x"6D6A6867",
									 -- x"69676667", x"67666768", x"68656260", x"5F5E5E5E", x"5C5C5E61", x"63646566", x"64656564", x"64686A6B",
									 -- x"6B6C6D6E", x"6E707375", x"797A7B7A", x"7B7F8080", x"8585878C", x"939DA6AD", x"A6A6A5A4", x"A09A9591",
									 -- x"95918D8F", x"92959FB0", x"BEBECACE", x"C2BEBFB7", x"B1ABBAB0", x"BBD1CEE9", x"F7F8F9F4", x"EFF1EFE5",
									 -- x"E4F0F6F7", x"F7E9DDE0", x"E3E3E5E7", x"E6E2DFDF", x"DAD8D6D6", x"D6D5D2CE", x"D1D1CDC9", x"C9CDD0D1",
									 -- x"D3D0D4D5", x"CFD0D4D1", x"D5D3D0CC", x"C6C0BDBB", x"BCBCC0C1", x"BDB5B3B7", x"B2B8BFC6", x"CCD0CDC8",
									 -- x"C9CDCAC1", x"B8B4B2B0", x"ABABAAA7", x"A39F9D9C", x"9A98938D", x"89858484", x"7C807A7B", x"79747975",
									 -- x"6E737269", x"6C736A6B", x"6B696165", x"6B68666A", x"66686968", x"625E5D5F", x"5D5A5955", x"4F4E5050",
									 -- x"4F4C4A4B", x"4B474341", x"41403C39", x"3A3D3830", x"302F2E2F", x"2F2E2C29", x"2C2A2725", x"24242322",
									 -- x"25221F1E", x"1F201F1E", x"21201E1E", x"1E1C1A18", x"191B1B1C", x"1B1C1D1F", x"1B1A1A19", x"19191A1A",
									 -- x"1C1C1A17", x"15161514", x"14151617", x"17171716", x"16161616", x"16161617", x"19181616", x"16161615",
									 -- x"14151413", x"14161513", x"13141414", x"13131414", x"13121214", x"13101012", x"0D0F1010", x"0F0E0E0E",
									 -- x"0C0B0C0D", x"0D0C0C0D", x"0D0E0E0E", x"0C0B0C0C", x"0D0D0D0E", x"0F100F0F", x"0D0C0C0C", x"0C0D0E0F",
									 -- x"0F0F0E0E", x"0F101111", x"10121211", x"1213120F", x"10121311", x"11131415", x"17161414", x"14151413",
									 -- x"15141312", x"11111112", x"15121112", x"110F0F10", x"12121313", x"14131314", x"13131313", x"14161819",
									 -- x"17181A1D", x"1E1E1D1D", x"20201F20", x"21232629", x"26232324", x"23202024", x"1D1F2123", x"24252424",
									 -- x"24282926", x"25282826", x"25282B2C", x"2B2A2C2E", x"2929292A", x"2F322F29", x"2C2E2F30", x"32353533",
									 -- x"D3D1CFCE", x"CECCCBCA", x"CBC5C4C5", x"C3C4C8C9", x"C8C9C9C9", x"C9C7C6C5", x"C4C2C0C1", x"C1BFBEBF",
									 -- x"C1C1C1BF", x"BEBFBFBD", x"BEBDBCBC", x"BDBDBAB8", x"B5B2B1B2", x"B3B3B3B3", x"B3B3B2B1", x"B1B2B3B4",
									 -- x"B2B1B1B0", x"ADAAABAD", x"ACAAAAAA", x"ACACABA9", x"A9A9A9A8", x"A7A7A8A8", x"ACAAA8A8", x"A9A8A5A2",
									 -- x"9A938C87", x"86878A8C", x"87847F7D", x"81878B8C", x"8D8C8885", x"85868583", x"7E7B7978", x"76736F6E",
									 -- x"706E6E6F", x"706F6F70", x"6C6B6968", x"68676767", x"6465676B", x"6C6C6C6C", x"6C6E6E6B", x"6A6C6F70",
									 -- x"73747574", x"74757779", x"7B7E8080", x"83888C8E", x"8D8D9299", x"9FA5ADB3", x"B1B2B6B9", x"B6ADA49F",
									 -- x"9B9C9A98", x"9797A3B5", x"C9CDDCDF", x"D4D0CFC6", x"BCB9B1BE", x"CDD5E9F4", x"FEFDF8EF", x"E7EAF1F2",
									 -- x"DCE6F9FF", x"F6E3DCDE", x"D9DADCDF", x"DEDBDADA", x"DBD8D4D1", x"D0CDCAC6", x"C7C8C8C7", x"C9CCCECE",
									 -- x"CECDD0D1", x"CECDCDCA", x"CECECECB", x"C5BFBAB8", x"B8B7BABD", x"BAB4B1B3", x"B4B8BDC1", x"C5C8C8C5",
									 -- x"C5C6C1B8", x"B0ADABA8", x"ABAAA8A4", x"A09D9C9C", x"96938F8B", x"87837E7B", x"756F786F", x"6876756C",
									 -- x"6A6B6766", x"73676B69", x"69646A6B", x"5F63636A", x"6C6E6A65", x"5B5B5D62", x"5C585755", x"5151524F",
									 -- x"4F4B4949", x"49464342", x"3D3F3E3A", x"37373632", x"32313030", x"302F2D2A", x"27272726", x"25252526",
									 -- x"26242121", x"21222121", x"22211F1E", x"1E1E1C1B", x"1B1C1C1D", x"1C1C1E1F", x"1C1C1C1C", x"1C1C1C1C",
									 -- x"16181A1A", x"19191714", x"17171818", x"18191919", x"17181819", x"19191818", x"19181818", x"17161515",
									 -- x"15161615", x"15161513", x"15151615", x"14131313", x"14131213", x"13111112", x"0E0F100F", x"0F0E0E0E",
									 -- x"0D0C0C0E", x"0E0C0C0D", x"0C0D0E0D", x"0C0B0C0C", x"0D0D0D0D", x"0E0F0F0F", x"0D0D0C0C", x"0D0E0E0F",
									 -- x"0F0F0E0F", x"10111111", x"12141413", x"14161715", x"10131413", x"12131414", x"18161515", x"15151413",
									 -- x"13121110", x"0F101112", x"110F0F10", x"11111113", x"12121313", x"14141415", x"16161616", x"16161617",
									 -- x"18191C1E", x"1F1F1F1E", x"20202020", x"21232527", x"22222223", x"22212122", x"1F202122", x"23222120",
									 -- x"22272926", x"24262726", x"26282B2B", x"2A2A2B2C", x"292C2E2D", x"2C2D2E2D", x"30313131", x"33353634",
									 -- x"DCD8D3D0", x"D0D1CECC", x"CDC6C3C2", x"C0C3C7C7", x"C9C9CACA", x"C9C7C5C4", x"C3C1C0C1", x"C1C0C0C0",
									 -- x"C1C1C0BE", x"BCBDBDBB", x"BEBBB9B9", x"BBBBB8B6", x"B0AEAEB0", x"B2B1B0B0", x"AFAEACAC", x"ADAEAEAD",
									 -- x"B1B1AFAD", x"ABACACAB", x"ADAAA9AA", x"ADAEACA9", x"A8A9A9A8", x"A7A6A7A9", x"ADABAAA9", x"AAA9A6A3",
									 -- x"9F99908A", x"8787888A", x"82817F7D", x"7C7D8184", x"8D8E8D8B", x"8784868A", x"827F7E7E", x"7D7A7979",
									 -- x"79777679", x"7B7A7978", x"75747372", x"71706D6C", x"6E6F7277", x"79787677", x"76787774", x"72737576",
									 -- x"7778797A", x"7A7B7E80", x"7F818384", x"868B9194", x"97979DA6", x"ACB0B7BF", x"BCBCC1C7", x"C3B7ACA9",
									 -- x"A8AAA8A5", x"A4A3ACBB", x"D9DFE8E5", x"D5CECABF", x"C1C8BFCB", x"D2DAF7FA", x"FBF7F1EC", x"EBF0FAFF",
									 -- x"E6DEE8F1", x"E4D9D8D7", x"D2D3D6D8", x"D6D4D5D7", x"D6D2CECC", x"CBCAC7C5", x"BFC1C1C1", x"C3C6C8C8",
									 -- x"C9CCCDCE", x"D0CDC7C6", x"C8CBCDCC", x"C7C0BAB7", x"B5B3B3B6", x"B7B3AFAE", x"B5B9BDBF", x"C1C2C2C1",
									 -- x"C3C1BBB1", x"ABA9A6A2", x"A4A3A19E", x"9C9B9B9C", x"96928D89", x"86807973", x"796D7277", x"6F676569",
									 -- x"6B626E5E", x"6169665F", x"60636860", x"65685E6A", x"60656468", x"63675F5B", x"5C585757", x"5453534E",
									 -- x"4F4C4947", x"46444241", x"3C3E3D39", x"36363432", x"3331302F", x"2F2E2C2A", x"25262827", x"25252729",
									 -- x"25232121", x"22222220", x"22211F1E", x"1E1E1E1D", x"1D1D1E1E", x"1D1E1E1F", x"1C1D1D1D", x"1D1D1D1D",
									 -- x"15181B1C", x"1C1C1A17", x"19191919", x"19191A1A", x"18191A1B", x"1B1A1919", x"18191A1A", x"18161616",
									 -- x"17181817", x"17171513", x"16161615", x"14141414", x"15141313", x"13121213", x"11100F0F", x"0F0F0F0E",
									 -- x"0E0D0D0E", x"0E0D0C0D", x"0C0D0E0E", x"0E0D0E0E", x"0E0D0C0C", x"0D0E0F0F", x"0D0D0D0E", x"0E0E0F0F",
									 -- x"0F0F0F10", x"11121211", x"12131312", x"12141616", x"11131413", x"13141413", x"15141413", x"13131212",
									 -- x"1211100F", x"0F101214", x"0F0E0E0F", x"11121314", x"12121313", x"13141515", x"15151617", x"18191919",
									 -- x"191A1D1F", x"21212120", x"20212121", x"21212223", x"1F202121", x"21232221", x"20212122", x"2221201F",
									 -- x"20262926", x"23242627", x"2728292A", x"2A2A2A2A", x"2B2D2F2E", x"2D2E2F30", x"31313130", x"32343432",
									 -- x"E4DFDAD6", x"D5D6D3CF", x"CFC8C4C3", x"C2C5C8C6", x"CACBCBCA", x"C9C6C4C3", x"C3C1C0C0", x"C1C0C0BF",
									 -- x"C1C1C0BD", x"BBBBBAB8", x"BDB9B6B5", x"B6B6B3B1", x"AEACACAE", x"AFAFAEAF", x"ACABABAA", x"AAAAAAA9",
									 -- x"AFB0AFAC", x"ADB0AFAC", x"ACABABAD", x"AFB0AEAB", x"A9AAABA9", x"A7A7A7A9", x"ACABAAA9", x"A9A7A4A2",
									 -- x"A39B938F", x"8C87878A", x"89888887", x"84808184", x"88898C8D", x"89868B92", x"8B888482", x"82828588",
									 -- x"85828285", x"88878583", x"7D7E7E7D", x"7C7A7774", x"78797D84", x"87868587", x"84858380", x"7F80807F",
									 -- x"7E7F8081", x"81828486", x"83858787", x"888C9297", x"9B999EA7", x"AEB2BBC4", x"C7C5C8CC", x"C7BCB4B4",
									 -- x"B8B6B1B0", x"B1B0B1B8", x"D4DCE4DF", x"D5D6D7D1", x"CDD2DED5", x"D7F1FBFB", x"FDF3E8E6", x"ECF2F9FF",
									 -- x"FFF0E5E0", x"D7D3D4D4", x"CFD0D2D3", x"D1CFD1D4", x"CECCC9C8", x"C7C7C5C3", x"C0BFBDBB", x"BBBDBFC1",
									 -- x"C4C9C8C9", x"CFCBC4C4", x"C4C8CCCB", x"C6C0BAB6", x"B7B1AFB2", x"B5B3AFAD", x"B3B7BCBE", x"BEBDBCBB",
									 -- x"BFBEB8B0", x"AAA7A3A0", x"9E9D9B99", x"97979797", x"958F8985", x"837F7872", x"706E6568", x"70686162",
									 -- x"5B61585C", x"55546E67", x"5E585F60", x"6262675D", x"686C6666", x"5E645C5A", x"5F5B5A58", x"5454534F",
									 -- x"4F4C4946", x"4442403F", x"3F3D3A38", x"38393530", x"3231302F", x"2E2D2C2B", x"28292928", x"27272727",
									 -- x"24232222", x"23232221", x"22212120", x"20202020", x"1E1F1F1F", x"1F1F1F1F", x"201F1F1F", x"1E1E1E1E",
									 -- x"1D1E1E1C", x"1C1D1D1C", x"1C1C1B1B", x"1B1B1C1C", x"191A1A1B", x"1B1A1A1A", x"181A1C1B", x"18171719",
									 -- x"18181818", x"18171513", x"15151615", x"15141515", x"15141314", x"15151413", x"1312100F", x"1011100F",
									 -- x"0F0D0E0F", x"0F0D0D0E", x"0E0F0F10", x"10101011", x"0F0D0C0B", x"0C0D0E0F", x"0D0D0E0E", x"0F0F0F0F",
									 -- x"10101111", x"12131211", x"10111111", x"10111213", x"13141413", x"12131412", x"14131313", x"12121111",
									 -- x"12111110", x"11121314", x"100F0F10", x"11121313", x"11121312", x"13151616", x"15151617", x"18181919",
									 -- x"191B1D20", x"22232424", x"21222221", x"201F1F1F", x"1E21211F", x"20242421", x"20202122", x"23232322",
									 -- x"21252726", x"24252627", x"27272829", x"2A2A2A2A", x"2D2C2B2C", x"3032312F", x"31313130", x"31333332",
									 -- x"E9E7E2DE", x"DCDBD7D3", x"D2CDCBCA", x"C8CBCDCA", x"CBCBCBCA", x"C8C6C3C2", x"C0C0BFBE", x"BEBEBDBC",
									 -- x"BFC0BFBD", x"BCBBB9B7", x"B9B6B2B0", x"B1B1AFAD", x"ADAAA8A9", x"ABABACAD", x"ABADAEAD", x"ABA9A9A9",
									 -- x"ACAEAEAD", x"AFB3B1AD", x"AAABAEB0", x"B1B0AFAD", x"AEAEAEAC", x"A9A7A7A7", x"AAAAA9A9", x"A9A7A5A3",
									 -- x"A0959194", x"938C8B92", x"95938F8C", x"8A898A8D", x"87878B8D", x"8C8B9096", x"96928F8D", x"8B8D9197",
									 -- x"95929295", x"98979492", x"85888A8A", x"8B8B8985", x"83838891", x"9595969A", x"98979594", x"94959390",
									 -- x"8E8F908E", x"8D8C8C8D", x"8B8C8E8F", x"9092989E", x"98969AA3", x"A9ADB4BB", x"C4C2C4C7", x"C4BDB9BB",
									 -- x"C0BFBBB8", x"B9B7B4B5", x"C6D0D8D6", x"D4DBE0DE", x"D5CDDCD0", x"D8F8F0EC", x"FFF8E5DD", x"E1E4E9F3",
									 -- x"FFFEECDA", x"D3CDCACD", x"CACACBCC", x"CAC9CCCF", x"CBC9C7C5", x"C4C1BEBC", x"C1BFBCBA", x"B9B8B9BB",
									 -- x"BDC2C1C3", x"C9C7C1C2", x"C1C5C8C5", x"C0BCB8B4", x"B7B1ADAF", x"B3B5B3B0", x"B0B3B7BA", x"B9B7B6B6",
									 -- x"B7B8B5AF", x"A8A3A09E", x"9D9C9A97", x"95939190", x"8C888482", x"827E7872", x"6D6F676C", x"65575F60",
									 -- x"5B60614B", x"7BBBBF90", x"A98D575D", x"5C566164", x"5D656565", x"5C5F5D5F", x"5E5B5B58", x"53525351",
									 -- x"4C4B4846", x"44434140", x"3F3D3A39", x"39393531", x"34333231", x"31302F2E", x"2E2C2A29", x"2A2A2826",
									 -- x"26262626", x"26252524", x"23232424", x"24232322", x"20202121", x"21212020", x"24232221", x"20202121",
									 -- x"2222201D", x"1C1E1E1D", x"1F1F1E1E", x"1E1E1E1F", x"1C1C1B1B", x"1A1B1B1C", x"1A1B1C1B", x"19181A1C",
									 -- x"18181819", x"19181615", x"15151515", x"14141415", x"13141516", x"17171514", x"15131110", x"11121110",
									 -- x"100E0F10", x"100E0E0F", x"0F0F1011", x"11121212", x"100E0C0C", x"0C0D0F0F", x"0D0E0E0F", x"0F0F0F0F",
									 -- x"12111112", x"13121111", x"0F0F1112", x"12121213", x"14151311", x"11131413", x"15151515", x"14131212",
									 -- x"11111212", x"12121212", x"11111111", x"12131312", x"12141413", x"14171716", x"19181615", x"14141415",
									 -- x"181A1C1F", x"22242626", x"24242423", x"211F1E1D", x"2122211E", x"20242523", x"20202122", x"23232424",
									 -- x"24252625", x"26272727", x"27272829", x"2A2B2B2B", x"2D2B2B2E", x"3132312F", x"32333231", x"33353635",
									 -- x"EAEAE6E2", x"E0DFDAD4", x"D1CECDCC", x"CACDCFCB", x"CBCBCAC8", x"C6C4C2C1", x"C0C0BFBD", x"BDBEBDBC",
									 -- x"BCBEBDBC", x"BBBBBAB9", x"B5B3AFAD", x"ADADADAD", x"ACA8A6A7", x"A8A9ABAD", x"ADAEAFAD", x"A9A7A7A9",
									 -- x"AAACADAE", x"B0B2B0AE", x"ABAEB1B4", x"B4B3B2B1", x"B5B4B2AF", x"ACA9A7A5", x"A7A7A7A8", x"A8A7A5A4",
									 -- x"9E959298", x"98919096", x"96979695", x"94959493", x"90909293", x"93939599", x"9B9A9A9A", x"98999DA2",
									 -- x"A3A1A1A3", x"A4A2A09E", x"93969898", x"999A9894", x"8F8F949E", x"A3A3A4A8", x"A9AAA9A9", x"A9A9A6A2",
									 -- x"9E9F9F9E", x"9D9B9C9D", x"9A9A9A9A", x"98989A9E", x"9B9A9DA3", x"A8ABADAE", x"B6B8BBBE", x"BEBBBBBC",
									 -- x"BBC0C1BE", x"BFBDBDC0", x"C2CACECC", x"CBCDCDCB", x"CDC4C6C5", x"CAD4D4D6", x"F1EFE3DA", x"DAD8DBE7",
									 -- x"EDEFDECE", x"D0CEC5C5", x"C5C3C3C5", x"C5C5C6C9", x"C6C5C4C3", x"C2C0BDBB", x"BDBCBBBC", x"BBB8B7B7",
									 -- x"BABDBEBF", x"C3C2C0C0", x"BFC3C4BF", x"BAB8B6B4", x"B5B0ABAD", x"B2B5B5B3", x"B3B3B4B5", x"B5B3B3B4",
									 -- x"B0B2B1AD", x"A7A19D9B", x"98979695", x"94918F8D", x"87868583", x"817C7671", x"73617575", x"6B776E61",
									 -- x"6A5A4D6D", x"A26F7C92", x"A7C19988", x"63656E4B", x"5C5D5F62", x"65625C56", x"5B595957", x"51515352",
									 -- x"4A4A4946", x"45454544", x"3D3F3F3C", x"38353536", x"34343433", x"33323130", x"312E2B2B", x"2D2D2B28",
									 -- x"28282827", x"27262625", x"22242525", x"24232323", x"23222323", x"24242322", x"24232221", x"21212121",
									 -- x"21222220", x"1F201F1E", x"1F1F1E1E", x"1E1E1E1E", x"1F1E1D1C", x"1C1D1E1F", x"1C1C1C1B", x"1A1A1B1D",
									 -- x"1817181A", x"1A191818", x"16161615", x"14131313", x"12141616", x"16161615", x"16141312", x"11111111",
									 -- x"100F0F11", x"100F0E0F", x"0F0F0F10", x"11121111", x"110F0D0D", x"0D0E0F10", x"0E0E0E0E", x"0F0F1010",
									 -- x"12121112", x"12121211", x"0E0D0E11", x"14141314", x"16151311", x"11141514", x"14151515", x"14131212",
									 -- x"10111213", x"13121110", x"10111212", x"13141412", x"12151615", x"15181816", x"17161514", x"13141415",
									 -- x"17181A1D", x"20232627", x"26272726", x"23211F1F", x"2322201F", x"21242524", x"20202021", x"21222324",
									 -- x"25252526", x"28292827", x"2728292A", x"2A2B2C2D", x"2B2D3031", x"2F2D2E31", x"31323231", x"33353634",
									 -- x"DEDEDAD8", x"DADBD6CE", x"CBCACAC8", x"C6C9CCC9", x"CAC9C8C6", x"C4C2C1C0", x"BFC0BFBD", x"BDBFBFBD",
									 -- x"BBBCBAB8", x"B7B8B8B7", x"B5B3B0AD", x"ABABADAE", x"AFABA9AA", x"ACAEAFB1", x"B2B1AFAC", x"A9A8A9AA",
									 -- x"ABABACAF", x"B0B0AFB0", x"AFB0B2B4", x"B6B6B5B4", x"B9B6B4B2", x"B0AEAAA7", x"A8A8A9A9", x"A9A8A6A4",
									 -- x"A19D9A9A", x"9A989798", x"969DA19F", x"9FA19F9B", x"9C9FA09E", x"9D9D9FA0", x"A0A1A3A5", x"A4A5A9AE",
									 -- x"ADABABAC", x"ABA9A7A6", x"A5A8A8A6", x"A6A8A6A1", x"9E9EA4AE", x"B2B0B0B4", x"B6B9BBBA", x"B8B7B4B1",
									 -- x"AEAFB0B0", x"AFAEAFB0", x"ACAAA9A8", x"A5A19FA1", x"A4A3A3A4", x"A9ADABA8", x"AEB3B7B9", x"B9BABBBA",
									 -- x"B6BCBDBC", x"BFC1C1C4", x"BEC4C5C5", x"C7C6C3C2", x"C4C2BDBF", x"BEB9BFC9", x"D0D7D2CE", x"D3D1D1DB",
									 -- x"DEDAD1CB", x"CCCEC9C4", x"C1BEBDBE", x"BFBFC0C1", x"BFBEBEBE", x"BDBDBCBC", x"B6B5B6B8", x"B9B7B6B7",
									 -- x"B9B9BCBE", x"BCBCBDBB", x"BCC0C0BA", x"B5B4B5B3", x"B1AEABAB", x"AFB2B2B1", x"B5B3B2B4", x"B3B1AFAF",
									 -- x"ADACABA8", x"A49E9996", x"91908F8E", x"8D8B8886", x"83838381", x"7D7A7877", x"7DB08E9C", x"81598A6C",
									 -- x"6E5C7C6C", x"373D796A", x"7D7494C6", x"C7ABBF8F", x"5F555450", x"5B575E5E", x"5B585958", x"53525351",
									 -- x"4C4D4B47", x"46474848", x"40414240", x"3B38383A", x"36363736", x"35333231", x"32302D2D", x"2E2F2E2C",
									 -- x"2A2A2A29", x"28272727", x"24252625", x"24242425", x"25252526", x"27272625", x"23242424", x"24242323",
									 -- x"23242523", x"23232220", x"1F1F1F1F", x"1E1E1E1D", x"20201F1E", x"1E1F1F1F", x"1E1E1D1C", x"1C1B1B1B",
									 -- x"1A18181A", x"1B1A191A", x"17171716", x"15141314", x"13161816", x"14141516", x"15151412", x"11101111",
									 -- x"11101011", x"110F0F10", x"100F0F10", x"12121211", x"12100F0E", x"0F0F1010", x"0E0E0E0E", x"0E0F0F10",
									 -- x"11111011", x"12131313", x"0F0D0C10", x"14151414", x"16161412", x"13161615", x"13141615", x"14121212",
									 -- x"11111213", x"13121111", x"0F111313", x"14141310", x"10141514", x"14161613", x"14141414", x"15161717",
									 -- x"1718181A", x"1D212426", x"26262726", x"24222121", x"23201F20", x"22232425", x"21212121", x"22232425",
									 -- x"24242527", x"28282829", x"282A2B2B", x"2A2B2D2F", x"2C2D3031", x"2E2C2F33", x"30313131", x"32353433",
									 -- x"CDCCC8C8", x"CED3CEC4", x"C8C7C7C5", x"C2C6CAC8", x"C9C8C6C4", x"C2C1C0C0", x"BCBDBDBB", x"BCBEBEBC",
									 -- x"BBBAB7B3", x"B2B3B4B3", x"B6B5B2AE", x"AAAAACAE", x"B3B0AEB0", x"B2B4B5B7", x"BBB7B2AE", x"ACADADAE",
									 -- x"AEACADB0", x"B0AEAFB2", x"B0AEAEB1", x"B4B6B5B3", x"B9B6B4B3", x"B3B2AEAA", x"ADAEAEAE", x"ACAAA8A6",
									 -- x"A2A3A09B", x"9C9F9F9C", x"A0A8A9A3", x"A2A8ABA8", x"A4A9AAA6", x"A4A6A8A8", x"A6A8AAAC", x"ADAEB4BA",
									 -- x"B3B2B2B2", x"B0ADABAC", x"AFB2B3B1", x"B2B5B4B0", x"ADADB3BD", x"C0BCBABD", x"BDC3C8C6", x"C2BEBDBC",
									 -- x"BEBFC0BF", x"BDBBBBBC", x"BAB8B6B6", x"B3AFACAC", x"AAA8A4A2", x"A6ADACA6", x"A8ADB0AD", x"ADB0B2B0",
									 -- x"B8B9B5B3", x"BABEBBB8", x"BBBEBDBE", x"C1C0BDBE", x"BBB9B8B3", x"B8BBB6BF", x"C1C6BEBA", x"C4C6C5CD",
									 -- x"D1CED3D1", x"C3BEC1BD", x"BDBAB7B8", x"B9B9B8B8", x"B9B8B7B6", x"B6B6B6B6", x"B2B0B0B2", x"B3B3B5B8",
									 -- x"B6B4B9BC", x"B6B6B8B5", x"B7BBBBB4", x"AFB0B1B0", x"AFADABAB", x"ACAEADAC", x"B2B0B1B3", x"B3AEA9A7",
									 -- x"AAA7A4A3", x"A09B9490", x"908D8A88", x"85817D7A", x"7A7A7A78", x"77797F83", x"8E774F71", x"87525186",
									 -- x"86847595", x"9EB4882C", x"435C6642", x"7E5494BE", x"A59E9E84", x"73525559", x"5E5A5A5A", x"5655544F",
									 -- x"50504D48", x"46484949", x"46444241", x"413F3C3A", x"3A3A3B3A", x"38363433", x"3332302F", x"2E2E2F2F",
									 -- x"2E2E2D2C", x"2B2A2A2A", x"292A2A29", x"2727282A", x"27262728", x"292A2827", x"2527292A", x"2B2A2827",
									 -- x"27282725", x"24252524", x"22222223", x"22212120", x"2020201F", x"1F1F1F1F", x"1F1F1E1E", x"1D1C1A19",
									 -- x"1C1A191B", x"1C1A1A1B", x"16171716", x"15151515", x"14181915", x"12121516", x"14141413", x"100F1011",
									 -- x"12101012", x"11100F10", x"11101011", x"13131211", x"1211100F", x"10101010", x"0E0E0D0D", x"0D0E1010",
									 -- x"10100F10", x"12131414", x"140F0D11", x"15161515", x"16161514", x"15181716", x"15161817", x"16141414",
									 -- x"12131313", x"13131313", x"10121313", x"1314110D", x"0D111311", x"1214130F", x"15161616", x"16161616",
									 -- x"18171718", x"1B1F2325", x"24242525", x"23222222", x"231F1E21", x"24232325", x"22212122", x"23252728",
									 -- x"23242627", x"2726282A", x"292B2D2C", x"2B2A2D2F", x"2F2C2B2E", x"30303133", x"31323333", x"34363533",
									 -- x"C9C5C2BC", x"BFC0BABD", x"BCBDBEBF", x"C2C6C6C5", x"C4C4C2BF", x"BFC1C0BD", x"C0BDBBBC", x"BEBEBCB9",
									 -- x"BBBDB8B3", x"B2B2B2B5", x"B6B3B1B1", x"B1AEACAB", x"AFB5BBBD", x"BDBEBFBF", x"BBBBBAB7", x"B5B3B2B1",
									 -- x"B3AEACAE", x"B0AEADAE", x"ACAFB0AF", x"AEAFAFAF", x"B6B4B3B4", x"B5B4AFAA", x"ABAEB1B3", x"B4B3ADA8",
									 -- x"A8A3A3AA", x"ADA8A5A5", x"A6ABADAB", x"AEB6B8B6", x"B6BABAB4", x"AFAEACA8", x"A6A9ABAC", x"B2BBBFBE",
									 -- x"BABAB9B7", x"B5B3B2B2", x"B6BCC4C9", x"C8C4C4C8", x"BEBDBFC4", x"C6C5C4C6", x"CAC9CDD2", x"D1CDCCD0",
									 -- x"CFCDCCCD", x"C4C0C7C2", x"C1C1BDB9", x"B5B4B0AC", x"A9ABABAA", x"A9AAA8A5", x"A7A7A9AB", x"ABAAABAE",
									 -- x"ACACAFB2", x"B3B2B3B6", x"B4B7B9B9", x"B9B9B5B1", x"B4B0B3BC", x"BCB4B1B6", x"B7B9B9B6", x"B3B5BCC2",
									 -- x"C8CACAC5", x"BFBAB9B9", x"BAB6B5B5", x"B0B0B4B5", x"B3B1B0B1", x"B1B0AFB0", x"ADACAEB0", x"B1B0B0B2",
									 -- x"B3B4B5B6", x"B4B2B1B1", x"B4B5B3B0", x"AFAFAEAB", x"A9AAA7A4", x"A5ABAEAD", x"AEB0B2B1", x"ADA8A5A3",
									 -- x"A29F9B96", x"9493908D", x"8D88877F", x"7F787976", x"6A7E7777", x"885B8876", x"3E3E6572", x"816A6C88",
									 -- x"5C706195", x"A1989780", x"456C6D5B", x"7D804593", x"93AE96C2", x"CDAB8769", x"515A5E5D", x"52565755",
									 -- x"57525255", x"464C494A", x"4B4C4A44", x"42444441", x"3D3C3C3B", x"3B3A3836", x"35353433", x"32313131",
									 -- x"3031312F", x"2D2C2E30", x"2E2C2C2C", x"2B29292A", x"2A2C2E2F", x"2F2D2B29", x"2B2A2A2B", x"2D2D2B28",
									 -- x"2A2A2A29", x"27262626", x"28262425", x"24222224", x"2221201F", x"1E1E2021", x"1D1C1C1C", x"1C1D1C1C",
									 -- x"191A1A1A", x"1A191817", x"17171615", x"171A1711", x"16171817", x"16141414", x"13131211", x"11111213",
									 -- x"0F101111", x"10101112", x"0F0F1114", x"17171512", x"12111210", x"0D10120F", x"0E0D0C0C", x"0C0C0C0C",
									 -- x"0E0F0F0E", x"0F131515", x"12131312", x"15181815", x"15141617", x"17151517", x"15161614", x"14151514",
									 -- x"0F101215", x"15131213", x"13131414", x"13121111", x"11131413", x"13151513", x"16161515", x"15161819",
									 -- x"18181717", x"191B1D1E", x"20202121", x"21212121", x"1F202021", x"21212020", x"24212124", x"25252628",
									 -- x"26262627", x"292A2A2A", x"2A2A2A2A", x"2C2D2D2D", x"302F2E2F", x"31323131", x"34353231", x"36383634",
									 -- x"CAC8C7BE", x"BCBAB4B9", x"BDBDBCBB", x"BCBEC0BF", x"BEBEBCB9", x"BABDBFBE", x"BEBDBCBC", x"BCBCBCBB",
									 -- x"B9BCB8B4", x"B5B4B2B3", x"B4B2B1B1", x"B0AEAFB1", x"B6BBBFC0", x"BEBDBDBC", x"BBBAB9B7", x"B6B5B4B3",
									 -- x"B4B0AEAE", x"AEAEAEAE", x"ADB0B0AE", x"ACADAEAD", x"AFAFB0B3", x"B6B6B4B1", x"B2B2B2B3", x"B6B9B7B4",
									 -- x"B0ABABB0", x"B2AFAFB3", x"B2B6B8B9", x"BCC2C5C5", x"C2C6C5BF", x"B9B6B3AF", x"ACAEADAC", x"B1BBC1C3",
									 -- x"C2C2C3C3", x"C2C1C1C0", x"C2C1C4CA", x"D0D3D5D8", x"D0CDCBCD", x"D1D3D4D5", x"D5D3D5DA", x"DDDFE5ED",
									 -- x"F2EBE5E2", x"D0C2C2BC", x"BEC0BEBA", x"B5B1ADA9", x"A9A8A4A0", x"9EA1A3A3", x"A8A7A7A6", x"A4A1A1A2",
									 -- x"A4A3A3A6", x"A9A9AAAC", x"AAADAFB0", x"B0B0AEAB", x"ABAAAEB7", x"B9B4B0B1", x"AEAEAEAD", x"AEB1B5B9",
									 -- x"BFC2C5C3", x"BEB8B5B3", x"B3B0B1B1", x"ADACAFAF", x"ADABAAAB", x"ACABABAD", x"ABA9AAAC", x"ADABACAD",
									 -- x"B1B1B2B3", x"B2B1B0AF", x"B2AFAEAE", x"AEAAA9AA", x"A4A5A4A1", x"A3AAADAC", x"AAAAA9A8", x"A6A3A09D",
									 -- x"97979694", x"92908B86", x"8B787F7F", x"747B7379", x"77A9A753", x"7A79706E", x"607D747F", x"90848774",
									 -- x"68887C8B", x"838591B2", x"9C717341", x"6B66492C", x"697B99A1", x"8DC1B884", x"78704E50", x"575A5859",
									 -- x"5B584E58", x"5B4F5949", x"524F4C4B", x"4745484E", x"45444241", x"403F3D3C", x"3A393736", x"36363738",
									 -- x"30323433", x"312F2F30", x"34333131", x"302E2D2E", x"2D2E3031", x"31302E2D", x"2D2D2E2E", x"2E2E2D2C",
									 -- x"2B2B2B2B", x"2A292928", x"29262526", x"25242325", x"24242323", x"22222222", x"1F1F1E1E", x"1E1E1D1C",
									 -- x"1C1C1B1B", x"1A191817", x"18181716", x"17181614", x"16171717", x"16151617", x"11121212", x"13131313",
									 -- x"11111212", x"11101112", x"12121214", x"17171614", x"14131412", x"0F111310", x"0F0F0E0E", x"0E0D0D0C",
									 -- x"0E10100F", x"10131514", x"12131312", x"13151513", x"18171717", x"15131213", x"14161614", x"13131210",
									 -- x"10101214", x"14131314", x"15141314", x"15151312", x"11131313", x"13151514", x"15151615", x"15161819",
									 -- x"19191919", x"1A1B1D1E", x"1E1E1F1F", x"1F1F1F1F", x"1E1F2021", x"22222222", x"211E1D1F", x"21222528",
									 -- x"29282829", x"292A2929", x"2B2B2A2B", x"2B2D2F30", x"2E2E2E2F", x"31323232", x"32343231", x"35363333",
									 -- x"CACCCCC3", x"BCB8B3B9", x"BDBEBEBC", x"BCBDBDBB", x"BCBBB8B6", x"B6B9BBBC", x"BABBBAB9", x"B7B6B7B8",
									 -- x"B7B9B6B3", x"B5B5B3B3", x"B4B3B2B1", x"B0AFB3B8", x"B9BEC1C1", x"BFBFBEBD", x"BBBAB9B8", x"B7B7B7B6",
									 -- x"B6B6B4B1", x"B0B1B1B0", x"ADAEAEAC", x"AAABABAB", x"ACADAFB2", x"B5B5B4B3", x"B5B5B4B4", x"B8BDBFBE",
									 -- x"B5B1AFB1", x"B0ADAEB3", x"B7B8BBBE", x"C2C6C9CA", x"C5C8C7C1", x"BCB8B4B0", x"B1B1AFAC", x"B0B9C0C2",
									 -- x"C0C1C2C3", x"C3C2C1C0", x"C1BEBDC0", x"C6CBCED0", x"D7DADBDA", x"DADCDFE0", x"DEDDDEE2", x"E6EBF4FC",
									 -- x"F4F5FAF8", x"DCC0BBB6", x"B9BCBDB9", x"B3ADA9A6", x"A2A29F9C", x"999A9A9B", x"9F9D9D9C", x"9A989899",
									 -- x"9C99989B", x"9EA0A1A2", x"A3A5A6A6", x"A7A8A7A6", x"A7A8ADB3", x"B7B5B0AB", x"A7A5A5A6", x"AAAEB0B1",
									 -- x"B7B9BBBC", x"B9B4AFAD", x"ADAAACAD", x"AAA8A9A8", x"A9A7A6A7", x"A7A7A7A8", x"A8A7A7A8", x"A8A7A8A9",
									 -- x"ADADADAD", x"ADADACAB", x"AFAAA9AD", x"ACA6A5A8", x"A1A2A19F", x"A1A5A7A6", x"A4A29F9D", x"9D9B9996",
									 -- x"93939290", x"8D89827C", x"7D7A7771", x"77678482", x"84AB7F72", x"80778284", x"757F6780", x"9C80756B",
									 -- x"8BAF8971", x"7091A3B3", x"9E8E4738", x"7338A46F", x"28527D7E", x"8895ACA6", x"A4AD957E", x"684E514F",
									 -- x"585D5C55", x"5557535A", x"53545351", x"4E4D4C4B", x"4D4B4846", x"46454442", x"41403E3C", x"3B3C3E3F",
									 -- x"37383938", x"35333333", x"37353435", x"34313132", x"31323334", x"34333231", x"30303130", x"2F2E2F30",
									 -- x"2E2E2E2E", x"2E2C2B2B", x"2C2A2929", x"28262626", x"25242424", x"25242321", x"22212020", x"201F1E1D",
									 -- x"1D1D1C1C", x"1B1A1918", x"1A191818", x"16151517", x"17171717", x"16161617", x"11121314", x"14131211",
									 -- x"12121212", x"11101112", x"13131314", x"16171615", x"16141513", x"10111310", x"0F101010", x"100F0F0E",
									 -- x"0F101110", x"11131413", x"14151615", x"14151615", x"17161516", x"14121214", x"11131312", x"11110F0D",
									 -- x"0F0F1113", x"13111113", x"13111011", x"14151311", x"12131413", x"14151514", x"15161616", x"16171819",
									 -- x"1A1A1A1A", x"1B1C1C1D", x"1C1D1D1E", x"1E1E1E1E", x"1F1F2021", x"21222222", x"201E1D1E", x"20222425",
									 -- x"25252627", x"292A2B2B", x"2B2C2C2B", x"2B2D3032", x"30303031", x"33343434", x"32363534", x"37363434",
									 -- x"CACCCFC7", x"C1BDB8BF", x"BABCBDBE", x"C0BFBCB7", x"B8B6B4B4", x"B7B9BABA", x"B8B8B7B5", x"B3B1B1B1",
									 -- x"B4B6B4B2", x"B6B7B5B5", x"B5B3B1B1", x"B0B0B3B6", x"BBBEC1C0", x"BFBFBEBD", x"B9BAB9B8", x"B7B7B8B9",
									 -- x"B7BAB9B4", x"B2B4B3B1", x"B0AFAEAC", x"ABABACAC", x"ABADB0B2", x"B3B3B3B3", x"B4B6B7B7", x"B9BEC1C3",
									 -- x"BCB7B3B2", x"B1AEAFB3", x"B4B3B6BC", x"C2C4C4C4", x"C7C9C8C4", x"C1BEBCB9", x"B7B8B7B5", x"B6BBBFC1",
									 -- x"C4C4C5C4", x"C4C2C0BE", x"BEBEBFBF", x"BEBFC2C5", x"CDD9E3E3", x"E0E1E3E4", x"E6E7E9EE", x"F2F5F9FC",
									 -- x"F5F4F8F8", x"DDC0BAB5", x"B4B5B5B3", x"AFAAA5A2", x"9D9C9A97", x"94939494", x"93929191", x"918F8F91",
									 -- x"92909092", x"94959799", x"9C9D9E9E", x"9FA0A1A2", x"A8ABAEAF", x"B0AFABA5", x"A3A1A0A2", x"A6ABACAD",
									 -- x"B3B2B1B1", x"B0ADABAA", x"A9A6A8AA", x"A7A6A6A5", x"A6A4A3A3", x"A3A1A1A1", x"A3A3A2A3", x"A3A3A4A5",
									 -- x"A8A7A6A6", x"A7A8A7A6", x"A9A5A5A8", x"A8A3A1A3", x"A3A3A19E", x"9EA0A09E", x"9F9D9996", x"95949392",
									 -- x"91918D88", x"84817C78", x"74717569", x"6D709A74", x"6F8B6773", x"75804C32", x"57768F61", x"76968392",
									 -- x"9AA98A7A", x"8591949B", x"83576F84", x"14276BC0", x"9C756860", x"7485A9D9", x"9E78BACD", x"BE939483",
									 -- x"6558585B", x"635A5A55", x"5654555A", x"5C5A5756", x"54514E4D", x"4D4C4A48", x"48474542", x"41414242",
									 -- x"41403E3B", x"38373839", x"36353536", x"36353536", x"35353636", x"36363535", x"33343434", x"33333333",
									 -- x"34343434", x"3432302F", x"312E2D2D", x"2D2B2929", x"27262525", x"26262321", x"23222121", x"21201F1E",
									 -- x"1D1D1D1C", x"1C1B1B1B", x"1D191718", x"17141518", x"19181716", x"15151515", x"13141414", x"13121110",
									 -- x"12121111", x"11111111", x"11111213", x"15161515", x"16131313", x"1011120F", x"0E0F1111", x"11101010",
									 -- x"10111212", x"12121212", x"12141616", x"15161719", x"14131313", x"13111214", x"0E0F0F10", x"10100F0E",
									 -- x"10101112", x"12101012", x"10100F10", x"12121211", x"13141414", x"14141413", x"16171717", x"17161718",
									 -- x"1919191A", x"1A1A1B1B", x"1C1D1D1E", x"1F1F1F1F", x"20202020", x"20202020", x"20202223", x"25242322",
									 -- x"21222425", x"2628292A", x"2B2C2E2D", x"2C2D3032", x"30303131", x"32333333", x"32363636", x"37363538",
									 -- x"CACBCDC7", x"C5C3BDC1", x"BAB9B8B9", x"BCBBB6AF", x"ADABABAF", x"B5B8B6B4", x"B5B4B2B1", x"B0AFAEAD",
									 -- x"AEB3B4B4", x"B8B9B7B7", x"B5B2B0B0", x"B1B1B1B3", x"BBBEBFBD", x"BBBAB9B7", x"B5B8B9B8", x"B5B4B6B9",
									 -- x"B6B9BAB6", x"B4B5B4B0", x"B5B3B1AF", x"AEADACAD", x"ABADAFB0", x"B1B1B2B3", x"B4B8B9B8", x"B7BCC3C7",
									 -- x"C1B9B1AF", x"AFAFB1B4", x"B3B2B6BE", x"C6C8C5C3", x"C7C8C7C5", x"C4C5C5C5", x"C5C5C4C2", x"C1C4C7C8",
									 -- x"C9C8C7C6", x"C5C3C0BE", x"BDBEBFBE", x"BDBEC0C1", x"C2CFDCE3", x"E6E8E8E7", x"E0E3E8ED", x"F2F4F3F0",
									 -- x"FFFAF4F1", x"DBC2BCB5", x"B0ADABAB", x"AAA7A29F", x"9F9B9590", x"8F8F9294", x"918E8C8B", x"89868484",
									 -- x"8686888A", x"8A898B8F", x"91929395", x"96989B9E", x"A5AAABA6", x"A3A4A29E", x"9E9D9C9D", x"A0A3A6A8",
									 -- x"ACA9A7A8", x"A8A7A6A7", x"A6A2A3A5", x"A2A2A3A2", x"9F9D9D9E", x"9E9B9A9A", x"9D9D9D9D", x"9D9E9FA0",
									 -- x"A4A3A2A2", x"A2A2A2A2", x"A2A2A2A1", x"A1A09E9C", x"A1A19F9D", x"9C9C9B99", x"9C9B9895", x"91909091",
									 -- x"8D8C8883", x"807E7B78", x"716B6F6E", x"66614D71", x"8C8D854A", x"5E451C1A", x"45807A79", x"766E7C85",
									 -- x"8891857C", x"8C8996A3", x"8B8BA2B8", x"83393D93", x"C69C8364", x"6460A0A5", x"7C7CC7AD", x"C4A4B6B7",
									 -- x"D29B7050", x"5A586463", x"655E5E66", x"645B5960", x"59575554", x"5453504D", x"4B4B4A48", x"47464545",
									 -- x"4443403E", x"3C3B3C3D", x"3A393A3C", x"3C3B3B3C", x"39393A3A", x"3A393838", x"3938383A", x"3B3B3937",
									 -- x"39393939", x"3A393735", x"33312F30", x"312F2E2D", x"2C2A2829", x"29292724", x"24232222", x"22212020",
									 -- x"1F1F1E1E", x"1D1D1C1C", x"1F1A1718", x"18161517", x"19181715", x"14141413", x"15141313", x"12111111",
									 -- x"11101010", x"11111111", x"0F101214", x"16161615", x"15121213", x"11121310", x"0F101212", x"11100F10",
									 -- x"11111212", x"12111010", x"0E0F1112", x"12121315", x"14121212", x"100F0F11", x"0E0E0E0E", x"0E0F1011",
									 -- x"13121213", x"12101012", x"0F101212", x"11111314", x"14141415", x"15151515", x"17181817", x"16161616",
									 -- x"17171818", x"18181818", x"1B1C1D1E", x"1E1F1F1F", x"2020201F", x"1F1E1E1E", x"21222324", x"25252322",
									 -- x"23242525", x"24242526", x"2A2C2F2F", x"2E2D2F31", x"2E2F2F30", x"31323333", x"31343434", x"3635353A",
									 -- x"CAC9C9C4", x"C5C3BBBD", x"BDBAB5B3", x"B4B4B1AC", x"A9A6A5A9", x"ACACA9A7", x"ACABAAAA", x"AAA9A7A5",
									 -- x"A5ACB0B2", x"B7B7B5B6", x"B5B3B1B3", x"B5B4B3B3", x"B4B6B7B6", x"B5B5B5B3", x"B0B3B5B4", x"B2B1B3B6",
									 -- x"B6B8B8B7", x"B6B6B4B2", x"B5B2B0AF", x"AEABAAAA", x"AEAEAEAE", x"ADADADAE", x"B2B5B4B0", x"AFB3BCC3",
									 -- x"C3BAAFAB", x"ABADAFB1", x"B1B4BAC2", x"C9CCCAC7", x"C5C5C4C4", x"C5C6C8C9", x"CECDCBC8", x"C7CACED2",
									 -- x"C8C6C4C2", x"C1C0BDBC", x"BEBDBBBA", x"BCBEBDBB", x"BCC0C8D3", x"DFE6E5E1", x"D7D9DBDF", x"E5E8E4DD",
									 -- x"E8ECF5F9", x"E0C3B9B0", x"ADA8A4A4", x"A5A39F9D", x"9F9A9594", x"93929190", x"8E8B8988", x"85817F7E",
									 -- x"7E808384", x"82818488", x"87888A8D", x"9093989C", x"A0A4A5A0", x"9C9D9E9C", x"9B9B9A9A", x"9B9DA0A2",
									 -- x"A2A0A0A3", x"A3A09FA0", x"A09B9C9D", x"9B9B9D9B", x"99979799", x"99979696", x"98999999", x"999B9C9B",
									 -- x"9E9E9E9E", x"9E9E9FA0", x"9FA1A09D", x"9D9E9D99", x"9A9A9999", x"999A9999", x"98999894", x"918F8F90",
									 -- x"8D8D8B86", x"817E7A77", x"70736C66", x"68533F73", x"7E817B81", x"3A232620", x"28667889", x"77817C89",
									 -- x"879AA274", x"838271A2", x"AA8D8F8F", x"A28C002C", x"71001345", x"5D7B8E9A", x"806ECCA3", x"8964898C",
									 -- x"94B57476", x"5D5C5E67", x"5D656A65", x"605F5D59", x"5B585656", x"5756524F", x"4C4C4C4C", x"4B4A4847",
									 -- x"42424242", x"41414040", x"40404042", x"42414041", x"3F3F4040", x"40403F3F", x"3F3E3D3F", x"41413E3B",
									 -- x"3B3A3A3B", x"3C3C3B39", x"36333234", x"35343232", x"2F2E2C2C", x"2C2B2927", x"26252524", x"24242322",
									 -- x"23232120", x"1F1E1D1D", x"1F1B1919", x"1A191817", x"17171515", x"15151413", x"13131211", x"11121314",
									 -- x"10101010", x"11121110", x"0F101315", x"16171716", x"17121316", x"14151513", x"12131413", x"110F0F10",
									 -- x"13121213", x"12100F0F", x"0E0E0F10", x"0F0F0F11", x"100F0F11", x"100F1012", x"12100F0F", x"0F0F1011",
									 -- x"11111112", x"110F0E10", x"0E101212", x"10101215", x"13131416", x"17171718", x"17181716", x"15151516",
									 -- x"16161717", x"17171717", x"191A1B1C", x"1D1E1E1E", x"1E1E1E1E", x"1E1F1F1F", x"21212020", x"21232423",
									 -- x"23242626", x"25252728", x"292B2D2E", x"2E2E2F30", x"2E2F3132", x"33343536", x"32353435", x"3736373C",
									 -- x"C6C4C4C0", x"C2C1B9BA", x"BCBAB6B2", x"B1B3B3B1", x"AEAAA7A6", x"A4A09E9D", x"A3A3A4A3", x"A19E9D9C",
									 -- x"9AA1A3A4", x"A8ACAEB3", x"B3B1B1B3", x"B3B2B1B2", x"ACAEAFAF", x"AFB1B1B0", x"ACADAFB0", x"B1B1B1B1",
									 -- x"B5B3B2B3", x"B4B2B1B1", x"B0AEACAD", x"ADABAAAA", x"AFAEACAA", x"A9A8A8A8", x"AEAEACA7", x"A5A8AEB2",
									 -- x"BCB7B1AE", x"AEAEAFB0", x"B1B9C1C5", x"C8CCCDCB", x"CAC9C8C7", x"C8C8C9C9", x"CCCAC8C6", x"C6C9D0D5",
									 -- x"D0CCC7C4", x"C1C0BDBC", x"BFBFBEBC", x"BCBDBBB8", x"B6B4B5BE", x"C8CECFCD", x"CECECDD0", x"D7DCD7CD",
									 -- x"C0CFE4EF", x"DBC3BAB0", x"ABA6A2A1", x"A09D9B9A", x"9A969395", x"95918A86", x"86848384", x"83807E7D",
									 -- x"7D7D7E7F", x"7E7E8185", x"82828588", x"8B8E9499", x"9A9D9F9D", x"9C9D9D9C", x"99989898", x"999A9B9C",
									 -- x"9D9A9A9C", x"9B969496", x"98939496", x"94949594", x"95939293", x"92919191", x"92939493", x"93959593",
									 -- x"95979A9A", x"98989A9D", x"9E9D9B9B", x"9B999897", x"94939293", x"94959696", x"95959493", x"918F8E8D",
									 -- x"8F8F8C86", x"817C7875", x"736E6E61", x"68718E69", x"786350AA", x"2024041C", x"1551798C", x"72758799",
									 -- x"C59B698B", x"8785B78F", x"8E9C4B70", x"8679613A", x"170A378C", x"4E908B5D", x"88A49195", x"8F6DBB8E",
									 -- x"A05902AC", x"A59B7754", x"5E64645E", x"6067655B", x"5D595655", x"5655514E", x"4E4F4F4F", x"4E4C4A49",
									 -- x"46454545", x"45454545", x"45444548", x"48474647", x"46464849", x"49494948", x"47464646", x"46464442",
									 -- x"41403F3F", x"40403F3D", x"3D3A383A", x"3B393634", x"31313131", x"302E2B2A", x"2B2A2929", x"28282726",
									 -- x"26252423", x"21202020", x"1D1E1E1C", x"1B1B1A19", x"18171616", x"16151413", x"12121110", x"10111314",
									 -- x"10101012", x"1312110F", x"0F111214", x"15151617", x"18131417", x"17161715", x"14151615", x"13121213",
									 -- x"14121212", x"110E0D0E", x"110F0E10", x"100F0E0F", x"0D0D0E11", x"11111214", x"14121112", x"11101012",
									 -- x"10101113", x"12100F10", x"10111111", x"10111214", x"15141517", x"18171719", x"17171615", x"14151617",
									 -- x"16161717", x"17181818", x"1818191B", x"1C1D1D1E", x"1E1E1E1E", x"1E1F2021", x"2122211F", x"20232423",
									 -- x"21232526", x"26282A2C", x"28292B2C", x"2E2F3030", x"30313233", x"33343536", x"34363537", x"3A38373C",
									 -- x"C1C0C0BD", x"C0C0B9BB", x"B5B7B7B4", x"B2B4B6B7", x"B3B0ABA7", x"A19C9C9F", x"A0A2A3A1", x"9C989697",
									 -- x"93979694", x"989FA7B0", x"ADADAEAE", x"ACA9AAAC", x"ABACACAB", x"AAABABA9", x"AAA9AAAD", x"B0B2B0AE",
									 -- x"B0ABA9AC", x"ADACACAD", x"ADABABAE", x"B0AFAEAF", x"ABA9A7A6", x"A7A8A9AA", x"ABABA8A4", x"A2A2A3A2",
									 -- x"A5A6A8AB", x"ACACABAC", x"B5C0C9C9", x"C8CBCFCF", x"CAC9C7C6", x"C5C4C3C2", x"C5C4C4C4", x"C4C8CFD4",
									 -- x"D7D1CAC4", x"C0BDBAB8", x"B4BBC0BE", x"B9B6B6B5", x"B1AEAEB2", x"B4B4B7BB", x"BDBCBCC0", x"CAD1CBC0",
									 -- x"C3C2C5CE", x"C9C3C1B5", x"AAA6A3A1", x"9E9A9898", x"98908A8B", x"8C89837F", x"807F7F81", x"817E7C7B",
									 -- x"7C7A797A", x"7B7C7E82", x"7F7F8184", x"86898E94", x"9497999B", x"9C9D9B99", x"95959495", x"97979796",
									 -- x"9D999797", x"938D8C8E", x"928E8F92", x"9190918E", x"928F8C8C", x"8B8A8A8B", x"8A8C8D8B", x"8B8D8C8A",
									 -- x"8E929595", x"9494979A", x"9B969497", x"97929194", x"91908F8F", x"90919191", x"92919191", x"92908D8B",
									 -- x"8A898680", x"7C7A7876", x"6E6B6A6D", x"7767687C", x"6D9F9D68", x"491C1418", x"0E2E718F", x"97889797",
									 -- x"868A8384", x"7F85655C", x"A485825E", x"817AB38A", x"158BC8A7", x"54669AB3", x"8F9B8D88", x"7B7189A5",
									 -- x"620065B7", x"45B2C09B", x"92725C61", x"665E595E", x"605C5856", x"57565350", x"52525251", x"4F4D4B4A",
									 -- x"4D4B4846", x"46474949", x"48484A4C", x"4D4D4D4E", x"4A4B4D4F", x"50505050", x"5050504E", x"4C4B4B4B",
									 -- x"4C494747", x"47464442", x"46423F3F", x"3F3C3836", x"34353737", x"35322F2E", x"302F2D2C", x"2C2B2928",
									 -- x"27262524", x"23232323", x"1C20221E", x"1C1C1C1B", x"1A181717", x"16151311", x"13121110", x"10111112",
									 -- x"11111213", x"1313100E", x"10101112", x"12131516", x"19131418", x"17171715", x"14161716", x"15151618",
									 -- x"14121112", x"100D0C0E", x"110E0D0F", x"100F0E0E", x"100F1012", x"11100F11", x"14131214", x"14111113",
									 -- x"12121417", x"16141314", x"14131313", x"13141515", x"18161618", x"18161617", x"16151514", x"14151618",
									 -- x"17171718", x"18191919", x"1818191B", x"1C1D1E1E", x"1E1E1E1E", x"1F1F2021", x"22242423", x"24252421",
									 -- x"22242627", x"2626282A", x"2828292A", x"2D2F3131", x"30313131", x"30303031", x"33353437", x"3A373539",
									 -- x"B5B4B4B5", x"B7B9B9B9", x"B5B3B1B1", x"B3B5B7B8", x"B8B6B0A6", x"9F9FA1A3", x"9FA0A1A1", x"9F9C9996",
									 -- x"94908F90", x"8F8E959F", x"A4A9ABAA", x"AAA7A4A6", x"A7A8A8A8", x"A9AAA9A6", x"A9A7A7A8", x"ABACACAA",
									 -- x"A7A5A5A7", x"A9A8A8A9", x"ABA9ABB0", x"B5B6B4B3", x"AEACAAA9", x"A7A5A4A6", x"A6A6A6A4", x"A1A0A1A3",
									 -- x"A4A09E9F", x"A3A5A4A2", x"ABB6C2C9", x"C9C7C6C7", x"C3C2C1C0", x"BEBCB9B7", x"B8B5B7BF", x"C4C7CED8",
									 -- x"D5D5D1C8", x"BFB7B3B2", x"B2B6B8BB", x"BCB6B1B3", x"B0AFAEAB", x"AAAAACAF", x"ADB3B5B6", x"B9BCBCBF",
									 -- x"C3C2C1CA", x"C8C2C1B2", x"A8A6A39F", x"9B989695", x"8F908686", x"857F8075", x"777C7A7D", x"75787475",
									 -- x"757B7D78", x"777B7C79", x"7C797B83", x"888A8B8E", x"90929391", x"91949696", x"94918F8F", x"90909294",
									 -- x"93908D8D", x"8D8B8A8B", x"89898989", x"88878686", x"82848686", x"86858484", x"85878787", x"8586898C",
									 -- x"8B8A8C8F", x"92919293", x"8F8F9091", x"91908E8D", x"8E8B898C", x"8D8C8B8C", x"8F898D8D", x"9288888A",
									 -- x"8882867F", x"76787877", x"6E72758D", x"7B5B407D", x"8D859E64", x"2A180600", x"0510596A", x"748C8E8E",
									 -- x"93A27478", x"807A7E73", x"5B4D9B84", x"9D7B9887", x"80746695", x"A15A7EB2", x"8B9488AA", x"4D397B3C",
									 -- x"04A7B8A3", x"537E90B6", x"769E7A58", x"63635F5E", x"5F5A5757", x"57555455", x"55505153", x"4F4E4F4E",
									 -- x"5050504F", x"4D4C4D4E", x"4E4E5052", x"52505255", x"50555857", x"56585754", x"59585553", x"53535353",
									 -- x"51504F4E", x"4C4A4949", x"48474542", x"42423F3B", x"393C3D39", x"35363737", x"302E2D2C", x"2D2C2B2A",
									 -- x"29292B2C", x"29232021", x"231D1D21", x"201F1E1B", x"1B1A1615", x"18181616", x"12151513", x"12121312",
									 -- x"10111213", x"13131211", x"14131112", x"13141413", x"16141416", x"17161516", x"16161616", x"16151515",
									 -- x"17151312", x"1111100F", x"10111111", x"0F0F0F10", x"11101111", x"12131212", x"12151514", x"14151512",
									 -- x"12121315", x"15131415", x"16151517", x"19181513", x"16161717", x"16161718", x"16161514", x"15161819",
									 -- x"17171718", x"1819191A", x"1C1C1B19", x"17181B1D", x"1E1E1E1F", x"20202020", x"22212123", x"25262523",
									 -- x"27262526", x"27282726", x"29282829", x"2A2B2D31", x"31323334", x"35353434", x"35373838", x"38373839",
									 -- x"AEAEAFB0", x"B1B2B1AF", x"B4B2B0B0", x"B2B4B5B6", x"B1B0ADA7", x"A3A1A09E", x"9FA0A0A0", x"9F9D9A99",
									 -- x"98908C8D", x"8D8B8E94", x"9CA2A6A8", x"AAA6A3A4", x"A6A6A5A5", x"A7AAA9A6", x"A6A5A3A3", x"A5A6A8A8",
									 -- x"A5A3A3A5", x"A7A7A9AB", x"A6A7A8A9", x"ADB1B1AD", x"A9ACADA9", x"A7A6A6A4", x"A29F9D9E", x"A1A2A09D",
									 -- x"9E9D9D9F", x"A1A29F9D", x"A3A9B1B6", x"B9BABBBD", x"C0BDB9B6", x"B4B4B4B4", x"AFAFB2B7", x"BEC5CDD2",
									 -- x"D7D3CCC0", x"B5AEABAA", x"B1B5B6B8", x"B9B4B0B3", x"AEACA9A6", x"A4A3A4A6", x"A8B0B3B4", x"B6B6B4B5",
									 -- x"BCB8B7C8", x"D1CBC6B9", x"ADA9A29D", x"99979796", x"888A8282", x"817D7E77", x"777C7D7D", x"7776777B",
									 -- x"7D7C7A7A", x"79777778", x"7A787A81", x"8788888A", x"898B8B8B", x"8C8E8E8C", x"8E8C8A8A", x"8B8A8B8C",
									 -- x"8D898686", x"85838282", x"81818181", x"81807F7E", x"7F7E7E7E", x"7F7F7F7F", x"7D7E7E7F", x"80828385",
									 -- x"8484868A", x"8C8C8C8D", x"8F8D8C8B", x"8B8B8A8A", x"89868586", x"88878787", x"8688868A", x"89868482",
									 -- x"83807971", x"76786C6A", x"6F5E849E", x"64375D3F", x"7B9C7B7C", x"596A4E2E", x"0D153A46", x"3F6A9183",
									 -- x"86704C89", x"798BA37C", x"93BCA1A2", x"A573948D", x"C8B8946F", x"78607490", x"7B898F9D", x"64061B17",
									 -- x"6184AFA9", x"537D7A5F", x"25A5C38A", x"58646366", x"605D5B5C", x"5C5A5959", x"5A565758", x"55535352",
									 -- x"52535353", x"53535455", x"53535659", x"5958595C", x"5A5E5F5D", x"5E616361", x"6462605F", x"5E5D5C5B",
									 -- x"58565657", x"55524F4F", x"4B4B4A48", x"46464544", x"43403B37", x"393C3B38", x"37353231", x"31323131",
									 -- x"2F2D2C2B", x"28252528", x"28222224", x"2221201D", x"1B1C1A18", x"19181618", x"14161614", x"13141413",
									 -- x"11111213", x"12121110", x"13131212", x"13141414", x"16151518", x"19171615", x"17161514", x"14141515",
									 -- x"17151413", x"1312100F", x"10111211", x"100F0E0E", x"10101011", x"12131312", x"13151616", x"16181817",
									 -- x"16151515", x"15131416", x"17171718", x"18181817", x"18191919", x"18171718", x"17161615", x"15161818",
									 -- x"18181818", x"1819191A", x"1C1C1B19", x"17181B1D", x"1F1E1D1D", x"1D1F2122", x"22212122", x"23242424",
									 -- x"25252526", x"28292929", x"2B2A292A", x"2A2A2C2E", x"31323334", x"35353536", x"36373737", x"3738393B",
									 -- x"AAAAAAAB", x"ACACACAB", x"ADABA9A8", x"AAACADAD", x"A8A8A6A4", x"A3A3A09D", x"A1A1A1A0", x"9F9D9C9B",
									 -- x"988F8A8D", x"908D8B8B", x"939A9FA2", x"A6A5A4A6", x"A9A9A9A9", x"ABACAAA7", x"A3A2A09E", x"9D9D9C9B",
									 -- x"A2A1A2A4", x"A4A4A5A7", x"A3A6A49F", x"A0A6A5A0", x"A0A7AAA5", x"A2A4A29E", x"A19E9C9E", x"A1A19E9B",
									 -- x"999A9B9D", x"9FA09F9E", x"A1A2A5AA", x"ADB0B1B2", x"B1B1B0AF", x"AFADABAA", x"AAACADAE", x"B4BDC1C1",
									 -- x"BBBBBAB6", x"B1ADAAAA", x"B0B3B3B4", x"B5B2B0B2", x"ACA9A5A2", x"A0A0A0A0", x"A3ACB0B1", x"B2B1AFB0",
									 -- x"B1B4B9CB", x"D5CDC9C9", x"B8B0A59B", x"9592918F", x"8687817F", x"7C777772", x"75777D7C", x"79747B83",
									 -- x"817A7980", x"80787477", x"7B797B81", x"86858485", x"85858686", x"88898784", x"88868585", x"84838284",
									 -- x"86838181", x"807E7C7C", x"7A7A7B7A", x"79787775", x"76757577", x"7A7B7977", x"75757577", x"7A7C7C7C",
									 -- x"7D7E8185", x"87868686", x"88878686", x"86878888", x"85838283", x"83828182", x"81897F86", x"7E80807B",
									 -- x"7B777876", x"746E6B77", x"6675899F", x"34569982", x"46888B74", x"84A38492", x"97361719", x"2D3796A2",
									 -- x"5C845E4C", x"80A28A75", x"A7A07D6B", x"7184866B", x"A1AEADA6", x"856E6810", x"3C7C94A9", x"B43169AB",
									 -- x"818BA3B5", x"5F779A8F", x"4F88A8B0", x"6F636766", x"64636363", x"63616060", x"5F5C5D5D", x"59585856",
									 -- x"55565758", x"5858595A", x"595B5E60", x"615F6061", x"63666664", x"666A6E6E", x"6D6C6A68", x"67656463",
									 -- x"635E5D5F", x"5E595758", x"54565550", x"4C4B4A4A", x"4B46403D", x"3F413F3B", x"3C393634", x"34353535",
									 -- x"33312E2C", x"2A28292B", x"2B252424", x"2221211D", x"1B1E1E1B", x"1A17161A", x"18181716", x"16171615",
									 -- x"13131313", x"13121110", x"12121313", x"13131415", x"16151719", x"1A181616", x"16151413", x"13151718",
									 -- x"16151414", x"14131110", x"10111313", x"12111010", x"11111112", x"13141414", x"13141515", x"16181817",
									 -- x"1B191817", x"15141417", x"1A1A1A19", x"18181A1B", x"1A1A1B1B", x"1A19191A", x"18181717", x"17171818",
									 -- x"19191919", x"19191A1A", x"1D1D1B19", x"17181B1E", x"1F1F1E1E", x"1F202122", x"22222222", x"22232526",
									 -- x"25252527", x"292A2A2A", x"2B2A2B2C", x"2B2A2B2D", x"30303031", x"33343536", x"36373737", x"37393B3C",
									 -- x"A3A2A1A1", x"A2A3A4A5", x"A5A5A4A4", x"A6A6A6A6", x"A6A5A39F", x"9EA0A09F", x"A1A1A1A0", x"9F9E9C9B",
									 -- x"97929196", x"98969392", x"989D9E9E", x"A1A2A3A8", x"A8ABACAB", x"AAA9A7A4", x"A2A09F9F", x"9E9B9691",
									 -- x"98999DA1", x"A2A1A2A3", x"A2A29F9B", x"9A9C9C9A", x"9DA0A19F", x"9E9F9D99", x"989A9D9D", x"9C9B9B9B",
									 -- x"9A9A9A9A", x"9A9C9EA0", x"9FA0A3A6", x"A8A8A7A6", x"A5A6A7A8", x"A9A9A7A6", x"ABABAAAC", x"B1B6B8B5",
									 -- x"B3B2B1B0", x"ADA9A7A7", x"ACAFAFAF", x"B2B0AEB0", x"ABA8A5A3", x"A4A4A5A4", x"A8AFB2B0", x"B0ADAAAB",
									 -- x"A5ADB3BE", x"C6C0BDC4", x"BAB1A499", x"928D8986", x"8484807C", x"77737270", x"72727A7A", x"7D768088",
									 -- x"86838893", x"948A8383", x"807F8084", x"87858281", x"83818081", x"8484807C", x"82818080", x"7E7C7C7E",
									 -- x"807D7C7D", x"7D7B7A7A", x"77787876", x"75747270", x"6E6E7074", x"79797570", x"71707071", x"73747575",
									 -- x"77787B7E", x"7F808081", x"80818283", x"84848382", x"8281807F", x"7E7D7C7C", x"7C847A80", x"7B7A7E78",
									 -- x"78737471", x"6E6C676B", x"6F614D56", x"694D0F66", x"848C687F", x"82A6BA80", x"A4C6846C", x"64142977",
									 -- x"99889571", x"74849285", x"98999F9E", x"83ACAF6A", x"8C928EA3", x"9628674E", x"2B828F8D", x"93407A75",
									 -- x"809790BF", x"9D6E8188", x"7B88909A", x"A9686E6A", x"6B6B6B6A", x"69676666", x"64616263", x"5F5E5D5A",
									 -- x"5C5C5C5D", x"5D5D5D5D", x"5F616364", x"63626364", x"68696A69", x"6A6E7070", x"72706E6D", x"6C6B6A6A",
									 -- x"6C646062", x"625E5D60", x"5D5E5C58", x"54525251", x"4D4C4A48", x"45444140", x"3F3C3937", x"37373635",
									 -- x"33323130", x"2D2B2929", x"2B262524", x"2222221F", x"1C201F1C", x"1B18171A", x"1A191717", x"17181715",
									 -- x"15151515", x"14141313", x"11121414", x"13131416", x"17161719", x"1A181616", x"15141414", x"1517191B",
									 -- x"16161514", x"14131312", x"11121314", x"14141414", x"13121213", x"14151515", x"14151516", x"16171717",
									 -- x"1B1A1918", x"17151517", x"1C1C1B1A", x"19191A1A", x"1A1B1C1C", x"1C1C1C1D", x"19191818", x"18181818",
									 -- x"1A1A1919", x"191A1A1A", x"1E1D1B19", x"18191C1E", x"1E1F2122", x"23222121", x"23242423", x"22232629",
									 -- x"27272728", x"29292A2A", x"2A2A2B2D", x"2C2B2C2E", x"2F2F2F30", x"31343637", x"35363738", x"393A3B3C",
									 -- x"9F9F9F9F", x"9F9FA0A1", x"A1A3A4A5", x"A5A5A4A5", x"A5A5A39E", x"9B9C9EA0", x"9FA0A1A1", x"A19F9E9C",
									 -- x"9C9A9B9E", x"9E9D9EA1", x"A7AAA8A4", x"A4A3A4A8", x"ABAFB1AE", x"ABAAAAAA", x"A29F9D9F", x"A19F9892",
									 -- x"9192969C", x"A0A2A5A8", x"A5A19F9E", x"9C9A9B9F", x"A19E9D9F", x"A09E9B9C", x"989B9FA0", x"9F9E9E9F",
									 -- x"9A9A9895", x"93939597", x"999C9FA1", x"A09F9F9F", x"A7A4A2A1", x"A2A6A9AB", x"AAA8A9AF", x"B5B7B7B7",
									 -- x"BBB5AFAB", x"A9A8AAAD", x"A7AAAAA9", x"ACACAAAB", x"AAA9A7A8", x"A9ABACAB", x"B1B6B7B3", x"B0AAA3A2",
									 -- x"A3A7A6A8", x"B3B6AFAF", x"ABA59C94", x"8F8A8581", x"7D7B7B77", x"74747375", x"73707879", x"7F7A8287",
									 -- x"868A949D", x"9E99928F", x"8A898889", x"8A878380", x"807C7979", x"7B7B7875", x"7A797878", x"7776787B",
									 -- x"78767577", x"77757373", x"72747573", x"7373716E", x"6A6A6B6F", x"73736F6A", x"6B6C6C6C", x"6B6B6E71",
									 -- x"6F717374", x"7677797A", x"7C7C7D7E", x"7E7D7B7A", x"7B7B7B7A", x"78777878", x"76787779", x"7B717773",
									 -- x"716B6B65", x"687A7D76", x"6E482A2B", x"36326A6E", x"774D1451", x"514A9A8D", x"6D98B9B7", x"C5CB5206",
									 -- x"70929591", x"A67A6689", x"6F848287", x"4D73867A", x"856E7F80", x"92B0A9C2", x"58406475", x"6E2F8477",
									 -- x"8D8F89A4", x"7B336788", x"99929399", x"9B746C6B", x"7372716F", x"6D6C6B6A", x"6A686A6A", x"66666662",
									 -- x"63636363", x"63636363", x"65666766", x"65666768", x"6A6C6D6D", x"6D6E6D6C", x"71727374", x"7472706E",
									 -- x"6E686667", x"67636264", x"6061605E", x"5D5E5D5B", x"5453514E", x"4B484544", x"43413E3C", x"3B3A3836",
									 -- x"34343332", x"302D2A28", x"2C282726", x"24252623", x"1F201E1C", x"1D1B1819", x"1C1A1818", x"19181716",
									 -- x"17171616", x"15151515", x"12131414", x"14141516", x"17171719", x"18171618", x"15151515", x"16171819",
									 -- x"17161514", x"14141515", x"13131313", x"14151616", x"14131313", x"14141414", x"16161617", x"18181819",
									 -- x"19181919", x"18161618", x"1B1A191A", x"1B1C1A19", x"191B1C1D", x"1D1D1D1D", x"1A1A1919", x"18181819",
									 -- x"1A1A1A1A", x"1A1A1B1B", x"1E1D1C1A", x"1A1B1D1F", x"1E1F2122", x"23222121", x"23242322", x"22232629",
									 -- x"28292929", x"29292A2A", x"2B2B2C2D", x"2D2C2C2E", x"2F2F2F30", x"32343638", x"34353739", x"3A3B3B3B",
									 -- x"9D9EA0A1", x"A09F9E9E", x"9C9FA2A2", x"A1A0A1A3", x"A0A3A5A3", x"A1A2A4A5", x"A2A3A4A6", x"A6A5A3A2",
									 -- x"A2A09F9F", x"9E9FA4A9", x"AEB2B2B1", x"B1AEADB1", x"BCBFC1BF", x"BDBEC0C2", x"B8B4B0B0", x"B1B0ABA6",
									 -- x"A19F9FA2", x"A6A9ADB0", x"B1ABA8A8", x"A49D9EA4", x"ABA5A4A9", x"AAA4A1A3", x"A3A3A3A4", x"A4A29F9C",
									 -- x"97979694", x"92919292", x"999CA0A1", x"A1A2A6A9", x"ACAAA9A8", x"A9AAACAD", x"ADAAABB2", x"B8B9B9BA",
									 -- x"B8B3AEAE", x"AEACACAE", x"A5A7A6A4", x"A7A7A4A5", x"AAAAAAAB", x"ACADADAD", x"AEB3B4B2", x"B0AAA19D",
									 -- x"9C9EA09B", x"A0A7A3A3", x"9F9B9590", x"8C86807C", x"7A767775", x"73757378", x"75727679", x"7F7E8285",
									 -- x"878E969B", x"9D9D9996", x"95928F8E", x"8C898481", x"7E797575", x"77767473", x"73727272", x"71717477",
									 -- x"74717172", x"72706D6C", x"6C6F7170", x"7071706D", x"6B6A6969", x"696A6969", x"66676867", x"6666696C",
									 -- x"6A6C6E6E", x"6F727576", x"75757474", x"75767777", x"74767775", x"73747576", x"73707672", x"756A6A6A",
									 -- x"676A6A7E", x"A6A68A8C", x"774A2004", x"00498B79", x"791D0012", x"22284367", x"744A408A", x"9497B7BC",
									 -- x"846A1448", x"730A3987", x"A077747C", x"7C9C828A", x"9FA98E8C", x"99948781", x"7E0D3443", x"43B2AF52",
									 -- x"6BA785A9", x"81588B86", x"C08198B5", x"9287787C", x"7A797674", x"7374726F", x"6F6E6F6F", x"6B6B6C68",
									 -- x"68676666", x"67686868", x"696B6B6A", x"696B6D6E", x"6D6E7071", x"716F6C69", x"6D6F7376", x"76746F6C",
									 -- x"6C6B6C6C", x"6B676565", x"64656563", x"63636260", x"5F58514F", x"504E4A47", x"4543403E", x"3D3B3937",
									 -- x"38373532", x"302F2E2B", x"2C292827", x"24262825", x"22221E1C", x"201F1A1A", x"1D1B1B1B", x"1B191818",
									 -- x"18181716", x"16161617", x"14151616", x"16161616", x"18171819", x"18161718", x"18171616", x"15161617",
									 -- x"17171716", x"16161718", x"17151413", x"14151515", x"15141313", x"13141414", x"16151517", x"1818191A",
									 -- x"1817181A", x"19171718", x"19181719", x"1C1D1B18", x"1A1B1C1D", x"1C1C1C1C", x"1B1A1919", x"18191919",
									 -- x"1A1A1A1A", x"1B1B1C1C", x"1E1D1C1C", x"1C1D1F1F", x"201F1F1F", x"1F202223", x"23232322", x"23242627",
									 -- x"27282929", x"292A2B2B", x"2D2D2D2E", x"2D2C2C2D", x"2D2E2E2F", x"30323334", x"33343639", x"3B3B3B3A",
									 -- x"9C9D9E9F", x"9E9FA0A1", x"A2A6AAA8", x"A5A5A9AE", x"ACB0B3B4", x"B4B5B4B2", x"AFAFAFAF", x"AEADACAB",
									 -- x"A6A3A1A2", x"A5A8AAAC", x"AFB5B7B9", x"BBBAB9BD", x"C9CDD1D2", x"D3D4D4D2", x"D3D1CFCF", x"CECDCAC7",
									 -- x"C3BEBABA", x"BBBBBBBC", x"C1BEBBB8", x"B3ADADB0", x"B8B8BABD", x"BBB5B1B2", x"AEAFAFAE", x"AAA5A2A0",
									 -- x"A2A09D9A", x"9999999A", x"9EA2A7AA", x"ADB1B6BB", x"B5B6B7B8", x"B8B6B4B1", x"B5B5B5B7", x"BBBFC0BF",
									 -- x"C1BDBBBD", x"BAB2AAA7", x"A7A9A5A1", x"A3A4A2A2", x"A7A9AAAB", x"ABAAAAAA", x"A8ABAAAA", x"ADABA4A1",
									 -- x"94929A97", x"949A9A9E", x"9D9A9691", x"8B847E7B", x"7D777975", x"7578747A", x"7A7B7A7F", x"8187898C",
									 -- x"94979CA1", x"A6A7A5A2", x"9B989490", x"8D8A8582", x"7F7A7778", x"7A797777", x"73737373", x"716F7073",
									 -- x"716F6F71", x"716F6C6B", x"6A6E706F", x"6F716F6B", x"6C6C6A68", x"6666696B", x"67686868", x"67666667",
									 -- x"65686B6A", x"6B6E7171", x"706F6E6F", x"70717272", x"6F737471", x"6F6F7172", x"706B7269", x"686D6A71",
									 -- x"766EB1DA", x"B4A5AA98", x"7E5F6156", x"3B60772A", x"3B18083B", x"2F16046A", x"46240D77", x"6A6C758C",
									 -- x"A4B28C19", x"07000858", x"797D7F8C", x"958B908F", x"8CC5AA93", x"64999016", x"1F8A5D3B", x"1B85601D",
									 -- x"268490CC", x"8995E881", x"7B6CAAA7", x"AA787B81", x"807F7D7B", x"7D7F7C77", x"75747573", x"6F70706C",
									 -- x"6D6B6969", x"6A6C6C6C", x"6A6D6E6C", x"6B6D6F6F", x"70707071", x"716F6C6A", x"6B6C6D6F", x"6F6D6A68",
									 -- x"6A6C6D6A", x"67676766", x"65676866", x"64626160", x"615B5553", x"524F4C4B", x"4643403E", x"3D3C3A39",
									 -- x"38383532", x"3132302D", x"2D2B2B29", x"25272824", x"2625201F", x"22221E1E", x"1F1E1F20", x"1E1B191A",
									 -- x"1C1B1A19", x"18181819", x"18181819", x"19191817", x"1818191A", x"19171719", x"1B1A1817", x"16171819",
									 -- x"17191A1A", x"19191919", x"19171616", x"16171716", x"17161515", x"16171717", x"17151517", x"1817181A",
									 -- x"19191919", x"18171719", x"18181819", x"1A1B1A18", x"18191B1C", x"1B1B1A1A", x"1B1A1918", x"18191A1B",
									 -- x"1A1A1A1B", x"1B1C1D1E", x"1D1D1D1E", x"1F202020", x"21201F1F", x"1F212324", x"24232324", x"25262726",
									 -- x"26272929", x"292A2B2C", x"2E2D2D2E", x"2D2C2C2E", x"2D2D2F30", x"31313131", x"34343638", x"3A3B3A39",
									 -- x"A5A5A4A3", x"A4A8ADB1", x"B4B8BBB8", x"B4B4BBC2", x"C6C8C9C8", x"C8C6C2BE", x"BCBBBAB8", x"B5B3B2B1",
									 -- x"A9A5A4AA", x"B2B5B3AF", x"B3B8BABB", x"BEBEBEC2", x"C6CBD2D8", x"DCDBD5CE", x"D1D4D7DA", x"DAD9D8D7",
									 -- x"DAD5D1D2", x"D2CFCBC8", x"CBCCCBC7", x"C2C1C2C3", x"C4CBD1D1", x"CCC6C2C0", x"BCC2C7C3", x"BBB5B6BA",
									 -- x"B7B2AAA4", x"A1A1A1A2", x"9FA4ABB2", x"B7BCC1C4", x"C2C1C0BF", x"BFBFBEBD", x"BBBFBFBD", x"C1CACECA",
									 -- x"CEC9C7C9", x"C7BFB8B5", x"ACADA7A1", x"A2A3A1A2", x"A5A7AAAA", x"A9A8A8A8", x"A9A9A4A2", x"A7A8A5A4",
									 -- x"A0939A9E", x"9FA6A2A2", x"9D9B9792", x"8C86827F", x"7E777A77", x"787C787F", x"81858288", x"87929599",
									 -- x"9A9A9DA6", x"ACADA9A7", x"9E9A9590", x"8D8A8682", x"807C7A7C", x"7D7C7B7B", x"79787877", x"736F6E70",
									 -- x"6F6D6E70", x"716F6D6C", x"6D717270", x"6F716F6B", x"6B6D6E6C", x"69686C6F", x"6B6B6B6B", x"6B696664",
									 -- x"5F636767", x"676A6C6C", x"71707070", x"6F6D6A68", x"6B6F706C", x"69696B6B", x"6A666A60", x"5E787684",
									 -- x"7E80898B", x"90979089", x"A1997670", x"878C7369", x"675B7883", x"666A501E", x"2A1E2C52", x"37526472",
									 -- x"76889987", x"51542201", x"276E5A78", x"8B8B8973", x"9A888D9B", x"9C9E771E", x"319DBD17", x"0527433C",
									 -- x"1C7F9690", x"8987C470", x"517EB8C4", x"A36D8384", x"84838282", x"8688847E", x"7B7A7A77", x"73747571",
									 -- x"73716E6D", x"6E6F7070", x"6A6D6E6C", x"6B6C6C6B", x"716F6E6F", x"6F6E6C6B", x"6D6B6967", x"67676868",
									 -- x"686B6A63", x"60636767", x"5F646766", x"62616262", x"5C5C5C5A", x"544D4B4D", x"4745413F", x"3E3E3D3C",
									 -- x"35363533", x"3333302C", x"3230302C", x"28292A26", x"28272321", x"24232122", x"20202223", x"201C1B1D",
									 -- x"201F1D1B", x"1A1A1B1B", x"1B1A1A1A", x"1B1B1A18", x"18181B1C", x"1B181718", x"1D1C1918", x"181A1C1E",
									 -- x"171A1C1D", x"1C1B1A1A", x"19191819", x"1A1A1A19", x"1A191818", x"191A1B1B", x"1B191819", x"1918191B",
									 -- x"1C1A1919", x"17161619", x"191A1A1A", x"18181818", x"1517191B", x"1B1B1B1B", x"1B1A1918", x"18191A1B",
									 -- x"1A1A1A1B", x"1C1D1E1E", x"1D1D1D1F", x"20212121", x"21212223", x"23242424", x"26252527", x"29292827",
									 -- x"27282929", x"29292A2C", x"2C2C2C2E", x"2E2D2E30", x"30313234", x"34343333", x"35353537", x"393A3A3A",
									 -- x"B0B1B5B9", x"B8B7BCC4", x"CAC9CBCD", x"CBC7C8CD", x"D6D3D1D2", x"D1CDC8C5", x"C0BEBEBF", x"BFBBB6B3",
									 -- x"B3B0AFB3", x"B7B9B9B9", x"BCBCBBBC", x"C1C4C3C0", x"C8CED4D5", x"D6DADBDA", x"D9DADAD9", x"D8D8D7D6",
									 -- x"D7D8D9D9", x"D7D6D6D7", x"D9D4CECC", x"CED1D3D3", x"CED0D2D1", x"CDC8C8CB", x"CDCECCCB", x"CDC9C6C9",
									 -- x"CAC6C3C1", x"BAAEA7A6", x"A7A8AFB3", x"B3B6BEC1", x"C5BFBBBA", x"BBBCBEC1", x"C0C1C1C3", x"C8CED1D1",
									 -- x"D0CFCBC9", x"CCCEC9C2", x"BAB8B0A8", x"A7ABA9A3", x"A6ADB4B6", x"B5B3B1AF", x"AAB1B3AE", x"ACAEADA9",
									 -- x"A3A6A9AC", x"AFB1AFAC", x"A6A5A197", x"8F898684", x"80848582", x"82888C8C", x"8C91979B", x"9D9FA2A4",
									 -- x"A7A3A2A5", x"ABACABA9", x"A29A9593", x"91908D86", x"82848583", x"81818283", x"878B8D8B", x"847D7A7A",
									 -- x"7E7A7675", x"7372706F", x"756B7179", x"6A716F6F", x"716C6D76", x"727D858A", x"94758386", x"8479898D",
									 -- x"93796C69", x"5D6A686B", x"6C686B6D", x"6B6B6567", x"67686969", x"69676665", x"65695B75", x"836C6883",
									 -- x"95837584", x"867B6C65", x"95766972", x"6B76668B", x"726D7A7D", x"7C699636", x"17090B04", x"1930186D",
									 -- x"48257361", x"85B89A75", x"2B0A296E", x"7183A392", x"8F6D609C", x"AE9E45A1", x"2A0692BE", x"680063AB",
									 -- x"7358AFCC", x"A7A98700", x"829DBAA1", x"75E99087", x"88858C87", x"8A8D9083", x"8284837C", x"78787876",
									 -- x"74727071", x"756C7673", x"726D7072", x"68706A6D", x"6A6C6D6E", x"69676862", x"62706563", x"65655964",
									 -- x"61636360", x"5E5F6265", x"5C606362", x"5D5A5B5E", x"58585753", x"504F4D4B", x"46403E40", x"413E3B3B",
									 -- x"3A373432", x"31303031", x"32312F2F", x"2F2E2B28", x"27272829", x"29272422", x"26232224", x"24221F1E",
									 -- x"1F202020", x"1F1F1E1E", x"1F1D1D1D", x"1D1D1A18", x"1B1B1B1C", x"1D1E1D1C", x"1C1A1A1B", x"1C1B1C1F",
									 -- x"1D1C1C1D", x"1D1C1D1F", x"1C1B1A1A", x"1B1D1C19", x"181A1A19", x"191B1B1A", x"18191A1A", x"1A191817",
									 -- x"1A18191B", x"1A171619", x"1B1B1A1A", x"1A1A1A1A", x"1C1D1E1D", x"1C1C1D1F", x"1A191919", x"19191A1A",
									 -- x"1C1B1B1D", x"1E1F1E1C", x"1E1F201F", x"1E1F2123", x"20222322", x"22232423", x"22252625", x"25272827",
									 -- x"28282929", x"2A2B2B2B", x"2F2C2B2E", x"30303031", x"32313234", x"33303032", x"3134383A", x"3B3C3B39",
									 -- x"C7C4C2C3", x"C2C1C5CA", x"D3D3D7DA", x"D9D5D6DA", x"DDDBDBDD", x"DDD8D2CE", x"CAC6C3C1", x"BFBCB8B6",
									 -- x"B8B5B3B4", x"B5B3B1B1", x"B9BEC2C2", x"C0C0C1C2", x"C6CCD2D4", x"D6DADAD8", x"D9DADAD8", x"D7D6D6D7",
									 -- x"D9D9DADB", x"DCDDDDDE", x"DEDAD6D4", x"D5D7D8D9", x"D6D7D8D7", x"D4D1CFCE", x"D4D9D6CF", x"D1D4D5D5",
									 -- x"DEDCDBDD", x"D9CBBBAF", x"AAA8AAAD", x"ADB1B8BA", x"BEBAB7B8", x"B9BBBDC0", x"C2C2C2C3", x"C7CBCDCC",
									 -- x"CFCDCAC9", x"C9C9C6C1", x"C3C2BDB7", x"B5B7B7B4", x"BABEC0BE", x"BCB9B7B5", x"B3BCC3C3", x"C2C3C3C1",
									 -- x"C5C4C3C2", x"C3C3BFBA", x"B5B1A9A0", x"98928E8D", x"8D929699", x"9DA3A4A1", x"A0A3A6A9", x"ABACAEAF",
									 -- x"ABA9A8AB", x"AEAEADAD", x"ACA5A19F", x"9C9A9790", x"8B8B8A88", x"888B9093", x"95959596", x"9795908C",
									 -- x"8A898681", x"7C777371", x"6E777368", x"76706D6C", x"67717D90", x"836F5576", x"66566C71", x"68778066",
									 -- x"8D7C7D90", x"755C6365", x"625A7263", x"67705F6E", x"68666361", x"5F606163", x"67597699", x"84839878",
									 -- x"887B6089", x"867F6870", x"717B7283", x"806E8A71", x"67656D63", x"69736178", x"8AA6901F", x"22251709",
									 -- x"020F2214", x"28795771", x"CC3A1014", x"2998A39E", x"938C77A8", x"BAB94BD3", x"6500ABB5", x"C16A1879",
									 -- x"9C875B8E", x"CD683E3B", x"82A17B95", x"8B91D673", x"76897E7E", x"86847C87", x"7E7E8081", x"807C7775",
									 -- x"7A727465", x"65656862", x"656A6561", x"69556866", x"676A6D63", x"67726066", x"63686263", x"5F615C61",
									 -- x"635D595C", x"60615F5D", x"5F5F5D5A", x"5857585A", x"57535152", x"514D4B4C", x"47454342", x"43423E3A",
									 -- x"39373533", x"32323232", x"32302E2E", x"2F2F2D2B", x"2A292928", x"28272524", x"25242425", x"25232223",
									 -- x"20202021", x"22222120", x"201F1E1E", x"1E1E1D1D", x"1D1E1F20", x"21212120", x"1F1D1D1E", x"1E1D1D1F",
									 -- x"1D1D1D1E", x"1E1D1E20", x"1C1D1D1C", x"1E1F1E1C", x"1C1E1E1D", x"1E1F1D1B", x"1D1D1E1E", x"1D1C1B1A",
									 -- x"1B1A1A1A", x"1918191A", x"1A1A1A1A", x"1B1C1C1D", x"1B1D1F1F", x"1E1C1B1B", x"1818191A", x"1B1C1D1D",
									 -- x"1E1D1D1D", x"1D1D1C1B", x"1E1E1F1F", x"1F202122", x"23242422", x"21222323", x"23252625", x"25272928",
									 -- x"2B2C2D2D", x"2E2E2D2D", x"312F2F31", x"31303031", x"32313031", x"31323538", x"3835363A", x"3B38393E",
									 -- x"D1CBC7C8", x"C8C7C7C9", x"D6D8DDE2", x"E3E0E1E4", x"E4E2E2E4", x"E4E1DCDA", x"D6D2CDCA", x"C6C2BEBD",
									 -- x"B8B6B4B4", x"B2B1B0B1", x"B1B9BFC0", x"BFC0C4C7", x"C6CCD2D5", x"DADEDDD9", x"D6D6D6D4", x"D1D0D1D3",
									 -- x"D5D5D6D9", x"DDE0E1E1", x"E4E3E1E0", x"E0E1E2E3", x"E2E4E4E2", x"E1E0DCD6", x"D9E2DED2", x"D3DDE1DF",
									 -- x"E6E6E7EA", x"E9DDC6B2", x"ADA6A4A6", x"A5A9AEB0", x"B3B1B0B2", x"B4B5B7B9", x"BBBDBFC2", x"C7CCCDCC",
									 -- x"CAC9C8C7", x"C6C4C2C3", x"C5C5C3C1", x"BFBFC0C1", x"C7C7C7C5", x"C4C6C7C7", x"C2CAD2D7", x"D6D5D7DA",
									 -- x"DBDBDBDC", x"DDDAD1C9", x"C3B9AEA8", x"A4A09E9F", x"A2A6AAAE", x"B3B7B5B1", x"B1B2B4B5", x"B6B7B6B6",
									 -- x"B3B2B3B5", x"B5B4B3B4", x"B5AFADAC", x"A7A4A19A", x"9B999693", x"9193979B", x"94939497", x"9B9C9996",
									 -- x"91929087", x"7F7A7672", x"746E7471", x"6D647073", x"7E816D71", x"7B61585A", x"62626355", x"6A67676D",
									 -- x"526E798D", x"7550605E", x"64626464", x"635A655F", x"63615E5B", x"5A5C5F62", x"59719074", x"6870677E",
									 -- x"81717791", x"8868706B", x"5E87406B", x"77958A79", x"6963505F", x"6578876E", x"6C8A5C71", x"2F050F1E",
									 -- x"7293A2BB", x"93674F04", x"33B7C13B", x"006C7575", x"898991A8", x"B1694EA6", x"626FE098", x"72A99F89",
									 -- x"7189896B", x"7C67C23E", x"7FA77E7C", x"ABB0CF85", x"59827B7B", x"747D7576", x"7876787D", x"7E777170",
									 -- x"716B7373", x"AE8E8B94", x"A0AFBBC0", x"9A96825D", x"5F69646A", x"69686363", x"605D6067", x"5C5B5C5F",
									 -- x"5E5B5A5D", x"5D5A5A5C", x"5D595654", x"54545453", x"554F4C4F", x"4F4A4749", x"43454441", x"40413D36",
									 -- x"38373634", x"34343433", x"32302D2D", x"2E2E2D2C", x"2D2C2A29", x"29292928", x"26262626", x"25242527",
									 -- x"21202021", x"2323211F", x"22222120", x"1F1E1F20", x"1E202222", x"22212223", x"22212122", x"21201F20",
									 -- x"20202022", x"22202122", x"1E202020", x"20222220", x"1F202020", x"21211F1B", x"20202121", x"21201F1F",
									 -- x"1D1D1D1B", x"1A1B1C1D", x"1B1A1B1B", x"1C1D1E1F", x"1D1E1F1E", x"1D1B1A1A", x"1C1D1D1E", x"1E1E1E1D",
									 -- x"1C1C1B1C", x"1D1E1F1F", x"1E1E1E1F", x"20222222", x"25262522", x"21232525", x"24262626", x"26282929",
									 -- x"2C2D2E2F", x"2F2F2D2D", x"2C2D2E30", x"302F2F30", x"30303133", x"33323233", x"39373739", x"39393B3E",
									 -- x"D3D0CFD1", x"D3D2D1D0", x"D6D8DDE2", x"E4E3E4E6", x"E8E5E3E4", x"E5E4E3E3", x"E0DDDBD9", x"D6D1CCCB",
									 -- x"C5C2BFBC", x"B7B3B3B5", x"B8BBBEBE", x"BDBFC1C1", x"C1C6CBD0", x"D5DAD9D4", x"CFD0D0CF", x"CBC9CACD",
									 -- x"CECFD1D4", x"D8DCE0E2", x"E7E8E9E8", x"E7E7E8E8", x"EAEDECEA", x"EBEDE7DE", x"DDE6E2D7", x"D7E0E4E4",
									 -- x"E4E5E5E4", x"E3DBC7B4", x"AEA6A3A3", x"A1A2A6A7", x"ABABABAD", x"AEAFB0B1", x"B3B6BABF", x"C5CBCCCB",
									 -- x"C4C3C4C5", x"C2BFC0C4", x"C2C1C1C2", x"C2C1C1C2", x"C5C4C3C4", x"C8CED2D3", x"D3D5DADE", x"DCDADCE0",
									 -- x"DCDEE0E3", x"E6E5E0DA", x"CFC0B2AD", x"ABA8A8AB", x"ACAEB0B1", x"B3B6B6B3", x"B4B5B6B8", x"B9B8B6B4",
									 -- x"B8B7B7B9", x"B9B7B6B6", x"B6B2B2B1", x"ABA7A49F", x"A3A19E9C", x"99969698", x"90949899", x"9897999B",
									 -- x"91938F87", x"817F7C78", x"70727275", x"73756C7E", x"82717F4F", x"61515D52", x"635C5F5D", x"5A535667",
									 -- x"5471666F", x"816B7066", x"64575D5D", x"595D635F", x"5C5C5C5A", x"5858595A", x"5B525B85", x"6A7D615B",
									 -- x"69877574", x"7D666A84", x"786C606B", x"8A5A55A1", x"6D6B6C62", x"71787161", x"A05A5792", x"72586593",
									 -- x"BD7D4A92", x"7990A88F", x"344E6EA4", x"76402048", x"49648DAD", x"5A6BE086", x"6BF2DE8E", x"46AED3B8",
									 -- x"CDBCC3A3", x"76FD867F", x"897C5480", x"A7B1880D", x"45786C6B", x"6F736871", x"73706F70", x"6F6B6867",
									 -- x"6B57559B", x"82ABC5D0", x"D5C2C7D2", x"CFB0D6BD", x"82635E59", x"5E656164", x"63626262", x"5E61615B",
									 -- x"585B5D5C", x"58565759", x"56545251", x"5252504E", x"534E4A4C", x"4C484544", x"4142413F", x"3E3F3B37",
									 -- x"39393836", x"36363534", x"3532302F", x"302F2E2C", x"2E2E2C2B", x"2B2D2D2C", x"2A292827", x"25252526",
									 -- x"24232323", x"2424211F", x"23242322", x"201F1F20", x"1F222424", x"22212223", x"24242425", x"24232221",
									 -- x"24242526", x"25232325", x"22232422", x"22232424", x"21212121", x"2324221F", x"21212222", x"22222221",
									 -- x"1E201F1D", x"1C1E1F1E", x"1D1D1C1C", x"1C1C1D1E", x"1E1E1C1B", x"1A1A1C1C", x"1F202020", x"201F1F1E",
									 -- x"1C1C1C1D", x"1E1F2021", x"1F1F1E20", x"22242423", x"25262624", x"24262828", x"27272727", x"27282A2B",
									 -- x"2C2D2E2F", x"2F2F2E2D", x"2C2E3133", x"32313233", x"30313334", x"34333333", x"32363835", x"363A3B39",
									 -- x"D9D8D9DB", x"DDDDDCDC", x"DBDDDFE2", x"E3E3E5E7", x"E9E6E4E5", x"E6E6E6E7", x"E7E5E4E4", x"E3E0DEDE",
									 -- x"DFDCD8D1", x"C7BCB6B5", x"B7BDC1C2", x"C0C0C1C1", x"C2C5C8CB", x"D1D5D3CE", x"C8C8C9CA", x"C8C6C7CA",
									 -- x"C8CBCFD1", x"D3D7DDE1", x"E6E8EAEB", x"EAE9E9EA", x"ECEEEDEB", x"EEF1ECE3", x"E3E9E7E1", x"E1E3E5E8",
									 -- x"E7EAE9E2", x"DCD5C8BA", x"ADA6A4A4", x"A09EA0A1", x"A4A5A7A8", x"A9AAAAAA", x"AFB2B5BA", x"BFC4C5C3",
									 -- x"C0BFBFC0", x"BDBABCC1", x"C0BEBEC1", x"C3C2C1C1", x"C1C0BFBF", x"C3C9CCCC", x"D7D5D7DA", x"DAD7D7DA",
									 -- x"DBDEE0E1", x"E3E5E6E5", x"DACAB9B0", x"ABA6A5A8", x"A4A7A9AA", x"ABADAFB0", x"AFB0B2B4", x"B5B4B2B0",
									 -- x"B5B3B3B5", x"B7B5B2B1", x"B2B0B1B0", x"AAA7A49F", x"9F9D9C9C", x"9A979697", x"92969A99", x"94929396",
									 -- x"90908D88", x"8685827D", x"79707A72", x"6D846A5A", x"7284635C", x"474D5F5D", x"5E675D5C", x"4C5F5B6D",
									 -- x"6A676970", x"875B5A55", x"4F665E57", x"575C5B58", x"56585957", x"55525151", x"56587F5B", x"7A967151",
									 -- x"41584633", x"5D616C6A", x"6B5A7470", x"7D7F848F", x"7A6C8178", x"796A7272", x"5042878C", x"A1A2A89D",
									 -- x"75639B84", x"929274B3", x"B245335C", x"48302050", x"1C245C2B", x"56C75859", x"A3C6C53B", x"A6D6C2AD",
									 -- x"8BA290B6", x"9F8975C0", x"B4946B53", x"57410005", x"867E6A67", x"635C656D", x"696A6762", x"5F5F5F5E",
									 -- x"527AA899", x"9EB0BAAF", x"A9A1B3B2", x"BDAC9FB4", x"C8C59D8D", x"89647363", x"5E58565C", x"655F5C61",
									 -- x"5C5E5C59", x"5A5C5954", x"55545251", x"50504E4D", x"504F4C48", x"494A4741", x"44414041", x"413E3C3C",
									 -- x"3B3C3B38", x"38393735", x"37353433", x"3433312E", x"2E2F2E2D", x"2D2F2F2C", x"2E2C2927", x"28282725",
									 -- x"27262626", x"26252322", x"21222323", x"21202021", x"22242625", x"23222324", x"24252526", x"26262524",
									 -- x"26262627", x"26242425", x"25262623", x"23242626", x"24232324", x"26272727", x"24232322", x"22222222",
									 -- x"1F212120", x"1F1F1F1E", x"1F1E1D1C", x"1B1C1C1D", x"1C1B1A1A", x"1B1C1E1E", x"1D1D1E1E", x"1F202121",
									 -- x"2221201F", x"1E1E1E1F", x"21202022", x"24262525", x"24262726", x"26282929", x"29292929", x"292A2B2D",
									 -- x"2E2E2F2F", x"30303131", x"2D2F3131", x"30303030", x"33333331", x"31323435", x"37393A39", x"38393B3C",
									 -- x"E4E3E3E2", x"E2E2E3E5", x"E5E4E4E3", x"E3E3E4E6", x"E6E4E5E7", x"E8E6E5E5", x"E8E6E5E5", x"E6E5E7E9",
									 -- x"E8E8E7E4", x"DBCEC5C2", x"BAC5CECD", x"C6C0C0C2", x"C4C6C7C7", x"CACFCECA", x"C3C1C2C5", x"C5C4C6C9",
									 -- x"C8CCCFD1", x"D1D5DBE1", x"E8EAEDEE", x"EDECECED", x"EDEEEEED", x"EFF1EDE7", x"E8EBEAE9", x"EAE7E6EB",
									 -- x"EAEDECE4", x"DAD1C6BC", x"ABA3A1A1", x"9C98999A", x"9B9EA0A0", x"A1A2A3A3", x"A8AAAEB2", x"B7BDBEBD",
									 -- x"BCBBBAB8", x"B6B4B5B7", x"B8B8B9BB", x"BEBFBEBC", x"BDBDBCBC", x"BEC1C1C0", x"C4C4C8CE", x"D2D3D3D5",
									 -- x"D8DDE2E3", x"E2E1DFDC", x"D9CCBEB4", x"ACA6A4A5", x"9EA1A4A5", x"A5A5A7A8", x"A7A8AAAC", x"ADADACAB",
									 -- x"AFADADB0", x"B2B0ACAA", x"ADABACAC", x"A8A6A4A0", x"9C999798", x"97949496", x"93929190", x"8F8C8987",
									 -- x"89888786", x"85827E7A", x"73787963", x"83886B75", x"70695880", x"8066436E", x"666E634C", x"5F62616D",
									 -- x"64665885", x"4C4A344E", x"32746B58", x"5A51524D", x"51535453", x"51515354", x"65543F56", x"61535992",
									 -- x"9062776D", x"65346679", x"6C6C659F", x"8398916D", x"5B767EA6", x"7B8E7F58", x"367B8D8A", x"86A5A28E",
									 -- x"818C5B85", x"8B818798", x"93641F3E", x"341A442D", x"1B242E3E", x"643D0F6B", x"8C6B5C15", x"223050B2",
									 -- x"A5ACA39D", x"897BD9B5", x"CAD1B685", x"6E644B79", x"6A5F5D58", x"645D5C57", x"595D5C56", x"52545553",
									 -- x"544C9CA3", x"AEB99F97", x"89A7B1B3", x"B3B4B6B3", x"A5C1C3B5", x"CEC4C0C9", x"BCB99B6A", x"58596366",
									 -- x"62646360", x"5F60605D", x"5A595652", x"4F4E4F50", x"4D4F4D48", x"484C4A43", x"48444245", x"433F3D3F",
									 -- x"3F403F3B", x"3A3C3A37", x"36353434", x"36353330", x"3031302E", x"2E2F2E2B", x"302E2B2A", x"2B2D2B28",
									 -- x"25252525", x"25242424", x"1F212223", x"22222222", x"22242525", x"23222223", x"22242626", x"26282726",
									 -- x"27262627", x"26242325", x"27282725", x"25272726", x"25242425", x"2626282A", x"28272624", x"23222222",
									 -- x"22212222", x"211F1E1F", x"1F1E1D1C", x"1C1D1E1F", x"191A1B1D", x"1F201F1E", x"1E1E1D1D", x"1D1E1F20",
									 -- x"22222222", x"21202121", x"23232425", x"26272727", x"25272827", x"26282827", x"2B2A2A2B", x"2B2B2C2F",
									 -- x"2E2E2E2F", x"2F303131", x"2F313231", x"32333434", x"2F323637", x"38393937", x"3B373639", x"38343840",
									 -- x"F0EFEEED", x"ECECEBEB", x"E9E8E6E4", x"E3E3E5E6", x"E5E5E5E7", x"E8E6E4E5", x"E6E5E5E6", x"E6E6E8EB",
									 -- x"E6E7E9EA", x"E7E1DCDB", x"D5DDE2DC", x"CFC5C1C0", x"C1C2C1BF", x"C2C7C8C7", x"C8C3C2C5", x"C7C7C9CC",
									 -- x"CFD1D4D5", x"D6D9DFE4", x"EBECEEEF", x"F0F0F0F0", x"F0F0F0EF", x"EEEDECEA", x"E9EBEAEB", x"ECEAE8EC",
									 -- x"EAEBEAE5", x"DDD4C8BF", x"AFA49E9E", x"9A969798", x"989B9C9B", x"9A9C9D9D", x"9FA1A4A9", x"AFB6B8B8",
									 -- x"B7B6B3AF", x"AEAEAEAD", x"ADB1B4B5", x"B7BBBBB9", x"BBBDBDBC", x"BDBEBDBB", x"B7B9BDC2", x"C5C8CBCD",
									 -- x"CFD4D9DB", x"DAD7D1CC", x"C9C5BDB6", x"AFAAA8A7", x"A1A2A2A2", x"A1A0A0A0", x"A1A2A3A3", x"A3A4A6A8",
									 -- x"A8A8A9AB", x"ABA8A5A4", x"A8A4A5A6", x"A4A4A49F", x"9F9B9898", x"96929092", x"93908D8D", x"8E8C8782",
									 -- x"817E7D7E", x"7D7A797B", x"806E7470", x"685E6667", x"48605C4B", x"744F5C55", x"745A7166", x"73636E5A",
									 -- x"6457454B", x"4C474A57", x"2A42825D", x"52594B55", x"4E505150", x"50515559", x"384B4942", x"64634135",
									 -- x"72728A8E", x"877E7A78", x"8A745D68", x"7C627B64", x"687D808E", x"7B6B9B4A", x"87918576", x"80A08C85",
									 -- x"9D4C3085", x"7B8C8A83", x"8D958B92", x"9261332B", x"2B1E182B", x"0A27584A", x"400C146E", x"AD1A2CBA",
									 -- x"BA8667B0", x"C281A0B1", x"A1ACAEAC", x"BDC08669", x"86937E48", x"58594F5F", x"5151504D", x"4C4C4D4D",
									 -- x"51458088", x"8CBA986B", x"88938CAF", x"7DADA5B4", x"B4BDB0B1", x"BEBEB9B7", x"C4BBC7CB", x"B8876A5C",
									 -- x"67646466", x"63606267", x"5E5C5956", x"53525151", x"4F504F4B", x"4B4C4B47", x"48474747", x"45434141",
									 -- x"4244423E", x"3D3F3E3A", x"38363435", x"36363432", x"33353330", x"2F31302D", x"30302E2C", x"2C2E2D2B",
									 -- x"26272726", x"24232426", x"23222223", x"24242423", x"22232324", x"24242323", x"22252626", x"27292928",
									 -- x"27262627", x"26252527", x"27282828", x"292A2926", x"26262727", x"26242629", x"29282625", x"24242424",
									 -- x"25212123", x"221D1D21", x"1F1F1D1D", x"1D1E1F20", x"1B1C1D20", x"22222120", x"22212120", x"201F1F1F",
									 -- x"21222324", x"23232425", x"24262728", x"28282829", x"282A2A28", x"27282928", x"2C2B2C2E", x"2E2D2D30",
									 -- x"2E2E2F30", x"30303030", x"35353433", x"34373837", x"34373733", x"2F2C2824", x"292C2D2D", x"2E33393C",
									 -- x"EFEFEFEF", x"F0EFEBE8", x"EAE9E7E5", x"E4E6E7E8", x"EAE8E7E8", x"E8E7E7E9", x"E6E7E9EB", x"EBE9E9EA",
									 -- x"ECEAEAEC", x"ECEBEAEB", x"E6E9E9E4", x"DED9D5D2", x"C5C6C5C3", x"C5CCCFCF", x"D2CBC7C9", x"CBCBCED1",
									 -- x"D8D9DADB", x"DEE2E6EA", x"EBEBEDEE", x"EFEFEFEF", x"F1F0EFEE", x"ECE9E8EA", x"E9ECEBEA", x"EDEDECED",
									 -- x"EDEBEAE8", x"E5DED2C8", x"B8A99F9E", x"9C9A9B9B", x"9B9D9E9B", x"9A9B9B9B", x"9C9EA0A3", x"AAB0B3B2",
									 -- x"B2B1ADA8", x"A9ACABA7", x"A8B0B5B5", x"B6BBBEBC", x"BDBFC0BF", x"BEBEBCBA", x"BDBEBFBC", x"BBBDC0C3",
									 -- x"C9C9C8C7", x"C9CBC9C7", x"BCBEBCB7", x"B1ADABA9", x"A6A29F9E", x"9E9E9E9D", x"A0A1A1A0", x"9FA0A4A7",
									 -- x"A2A3A6A7", x"A5A19F9F", x"A39F9FA1", x"A0A2A29E", x"A09C9A9B", x"99938F90", x"8D8C8B8B", x"8A888481",
									 -- x"807B787A", x"79777B83", x"78687086", x"63678068", x"525D4C65", x"6060565D", x"5A515459", x"5B5D5653",
									 -- x"2C3B182E", x"4D4B3448", x"38218370", x"4D48554C", x"4E4F504F", x"4D4D5053", x"2F4A4C43", x"62596044",
									 -- x"312B565B", x"5C648091", x"8B9B9787", x"7E756665", x"767D7578", x"9BA43F86", x"81698391", x"9A667E86",
									 -- x"5D3EAF95", x"777A888C", x"977A8684", x"73A7B889", x"81745D6F", x"5F2C133D", x"24503D93", x"C08116B9",
									 -- x"884396A1", x"692F6CA0", x"9598B4AE", x"BEA2AED1", x"CAB3BF86", x"4A4E5D4D", x"524C494B", x"4C4A4A4D",
									 -- x"41516866", x"898F8C89", x"7E8D726F", x"52606856", x"8E7F9DB0", x"98AFB2C8", x"C5BFB9A3", x"B0D1CC90",
									 -- x"6C5D5761", x"67636064", x"5E5D5B5A", x"59575350", x"5351504F", x"4D4A494A", x"474A4B49", x"484A4843",
									 -- x"45464540", x"4042413D", x"3E3B3838", x"38393736", x"36373632", x"32353531", x"2F31302D", x"2B2C2C2B",
									 -- x"2B2C2C29", x"26252629", x"27262423", x"24242423", x"24242526", x"27272726", x"23252626", x"27292A28",
									 -- x"27262627", x"2726282A", x"2627292A", x"2D2D2A25", x"29292B2C", x"29252629", x"27262524", x"24252627",
									 -- x"27212024", x"221B1C22", x"21201F1E", x"1D1E2021", x"201F1E20", x"21232322", x"21222323", x"24242423",
									 -- x"23252626", x"24232424", x"2527292A", x"2928292A", x"2B2C2B29", x"282A2B2B", x"2D2C2D2F", x"2F2D2E30",
									 -- x"30313233", x"33333231", x"32312D29", x"282A2926", x"262B323B", x"4B60717A", x"7A8C928A", x"8EA1A79F",
									 -- x"EEEEEEEE", x"EDECEAE9", x"EAE9E8E8", x"E8E8E7E6", x"E7E8E8E8", x"E8E7E7E7", x"E6E7E9EC", x"ECEAE9E9",
									 -- x"E9EAEAEB", x"ECEDEEEF", x"EBEDEDEA", x"E6E4E6E9", x"DAD6D3D3", x"D5D6D8DA", x"DAD5D1D0", x"D1D3D9DF",
									 -- x"E1E3E5E7", x"E9EAEAEA", x"EDEEEEEE", x"EFEFEFF0", x"EDEDEDED", x"ECEBE9E9", x"EAE9E9EB", x"EEF0F0EE",
									 -- x"EFEFEDEB", x"E8E4DDD7", x"C8B7A7A3", x"A5A4A2A1", x"A1A0A09E", x"9D9C9B9A", x"9BA1A5A6", x"A7AAACAC",
									 -- x"A9ACACA9", x"A9ACABA9", x"A8AEB5B9", x"BCBFC0BF", x"C1C3C1BB", x"B8BABDBD", x"BEBFBFBD", x"BBBBBEC1",
									 -- x"C4C7C7C4", x"C3C5C5C2", x"BBBAB6B2", x"B0AFACA9", x"A4A19E9D", x"9F9F9E9D", x"9FA1A19E", x"9FA09B94",
									 -- x"9D9FA1A0", x"9FA0A09F", x"A2A2A2A2", x"A2A1A09F", x"A49D9EA2", x"A09A9590", x"8E8A8984", x"84877F7B",
									 -- x"7880777A", x"74777672", x"7A37656A", x"67655853", x"5958515F", x"635A5354", x"846F5855", x"5358583C",
									 -- x"26221705", x"00050A26", x"15287F7A", x"897B4C45", x"52534658", x"4D495932", x"275E503B", x"595B294F",
									 -- x"21271E2E", x"4E544355", x"72797E75", x"7C758198", x"80827B6F", x"6A805878", x"6C748274", x"737C6E5E",
									 -- x"30638098", x"507F8698", x"928B8381", x"9592A291", x"96B0B197", x"C2AD4E4C", x"30050FB8", x"B6741CC1",
									 -- x"4D84CC3B", x"0F81334C", x"8A8895B7", x"928E7A9C", x"B4C2BED2", x"76373A3C", x"3F4C484B", x"40353A40",
									 -- x"423E606D", x"7E617DA0", x"BCACA27C", x"899FC09C", x"875BA0A9", x"A19FA8A7", x"97978C6D", x"779BB9AE",
									 -- x"C3BC8858", x"5C625F63", x"6159585B", x"57555654", x"5252504B", x"4C504F4C", x"484D4A45", x"484B4643",
									 -- x"4A474443", x"43444342", x"3D3D3D3C", x"3B393938", x"34343638", x"38353434", x"34333231", x"302F2D2C",
									 -- x"2C2C2B2A", x"29282726", x"28282726", x"25252627", x"26252425", x"26272625", x"26272727", x"292B2C2B",
									 -- x"2A292726", x"26272727", x"272A2C2A", x"292B2A26", x"292B2B29", x"27282826", x"26242426", x"26242426",
									 -- x"24222122", x"22211F1F", x"20212120", x"1E1C1C1C", x"1F1F2020", x"21222324", x"24232426", x"26252425",
									 -- x"25262728", x"29292928", x"2B2B2C2D", x"2D2B2A29", x"2B2C2C2C", x"2A292A2B", x"2B2D2F2B", x"30303632",
									 -- x"30313236", x"3234282D", x"2D2F5D71", x"7C6D627B", x"8E8FA4B5", x"B3AAB8A7", x"B9AFB1B6", x"BAB3A19C",
									 -- x"EFEFEEED", x"EDECEBEB", x"EAEAE9EA", x"EBECECEB", x"E9EAEAE9", x"E8E8E8E8", x"E7E7E8EA", x"E9E8E8EA",
									 -- x"E9EAEAEB", x"EBEBEDEE", x"EDEEEFED", x"EBEAEBED", x"E7E3E1E1", x"E1E0E0E1", x"E3E2E2E3", x"E2E1E3E7",
									 -- x"E7E8EAEB", x"ECEDEDED", x"EDEEEFEF", x"F0EFEFEF", x"EDEDEDED", x"EDEDEDED", x"EDEDEDEE", x"F0F1F1F0",
									 -- x"EEEEEDEB", x"EAE8E2DD", x"D5C5B5AE", x"AEADACAD", x"A7A7A8A9", x"A8A7A5A4", x"A5A9ACAD", x"AEB0B0AF",
									 -- x"B2B0ADAC", x"ABAAABAC", x"ADB3B9BD", x"C1C3C4C2", x"C3C4C2BE", x"BBBBBDBF", x"C1C0BEBD", x"BDBEBFC0",
									 -- x"C2C6C9C7", x"C5C5C2BD", x"BFBCB8B5", x"B3B1AFAD", x"A9A5A1A0", x"A1A3A4A5", x"A1A0A0A0", x"A09F9F9F",
									 -- x"989B9F9F", x"9E9EA0A3", x"A1A1A1A1", x"A1A09F9E", x"9C9EA3A3", x"A09F9C95", x"8B878883", x"82837B7A",
									 -- x"7A767873", x"75727384", x"4D435949", x"66473F4E", x"52666F5A", x"7A5A464B", x"54385233", x"4043380D",
									 -- x"06010201", x"1B39593C", x"1742856D", x"75896E86", x"5B46574F", x"5654583E", x"42634B47", x"564F6874",
									 -- x"6F403C3B", x"3B332F26", x"3A557888", x"66737572", x"66705A70", x"7379717E", x"5D6F7B85", x"9081624C",
									 -- x"2C5D7293", x"4E7D9176", x"79889A8F", x"93798FA5", x"A19D99A2", x"A5BDDBCA", x"BA87103A", x"E2A372A2",
									 -- x"67A99151", x"CE9B7646", x"5D668C9A", x"7C75758E", x"AEB2B2C7", x"A27F7A73", x"6E4A3F4A", x"6F82843D",
									 -- x"33483D62", x"75638188", x"A286927B", x"7E879CCF", x"9D919E98", x"AB7795A2", x"7588669F", x"9D7DA2A4",
									 -- x"ABBFC9C1", x"774A5E61", x"5A595B5A", x"54555854", x"5B535052", x"524E4E53", x"584E494E", x"514B484F",
									 -- x"4D4C4A49", x"49484745", x"41403F3D", x"3B3B3C3C", x"3B393939", x"39373637", x"35333130", x"2F2F2E2E",
									 -- x"2C2B2B2A", x"2A292929", x"2A2A2928", x"26262627", x"29272627", x"28292827", x"26262726", x"282B2B2A",
									 -- x"2C2A2928", x"29292A2A", x"272A2B2A", x"2A2D2C29", x"2A2B2B29", x"28292928", x"25242426", x"27262628",
									 -- x"26242324", x"23212020", x"20212323", x"22212121", x"21212121", x"22232425", x"25242527", x"27262627",
									 -- x"29282828", x"28292B2B", x"25272A2D", x"2E2E2D2C", x"2B2A2C2B", x"2B2C2A2B", x"30242C37", x"2F342725",
									 -- x"2D424838", x"3A44536D", x"8089AC98", x"9CB6BDA5", x"AEB1A0A2", x"A7A2A3AC", x"B1B0B0AF", x"ADA8A09B",
									 -- x"F0EFEEED", x"EDEDEDED", x"ECEBEBEC", x"EEEFEFEF", x"EBEBEBEA", x"E9E8E8E9", x"E8E7E7E8", x"E8E7E9EB",
									 -- x"E9EAEAEA", x"EAEAEBEC", x"ECEDEDED", x"ECEBECEC", x"EDEBEAEB", x"EBE9E8E8", x"EBECEFF0", x"EEEBEBED",
									 -- x"EBEBECED", x"EEEEEDED", x"EDEEEFF0", x"F0F0EFEE", x"EEEEEDED", x"EDEEEFF0", x"EFF0F0F0", x"F0F0F0F1",
									 -- x"EEEFEEEC", x"ECEBE8E4", x"E0D5C9C3", x"BFBBBABB", x"B9BABBBB", x"B9B7B4B1", x"B2B4B7B8", x"BBBDBDBB",
									 -- x"BDB8B6B7", x"B6B2B1B4", x"B4B9BEC2", x"C4C6C6C5", x"C7C6C5C5", x"C3C2C3C6", x"C8C4BFBD", x"BDBCBBB9",
									 -- x"BBC0C4C4", x"C3C4C1BE", x"BFBBB7B7", x"B6B3B2B4", x"B6B3ADA8", x"A6A5A5A5", x"A6A3A3A6", x"A39E9DA1",
									 -- x"9B9DA2A6", x"A5A3A6AC", x"A7A7A8A8", x"A7A5A4A3", x"9BA4ABA6", x"A1A4A297", x"908B8C88", x"86847D7E",
									 -- x"80736D6D", x"6E6B724C", x"60443330", x"24241D2D", x"3A1B282D", x"5E3D3546", x"50495E49", x"5D853222",
									 -- x"25222F47", x"6E8F8790", x"53505C6A", x"987F7B6D", x"8A704A52", x"4F545C3E", x"1B3F594D", x"5A4A5770",
									 -- x"523E3530", x"313A0A30", x"37534069", x"66686B60", x"25548490", x"A36A5E91", x"797A8A88", x"707B4B6B",
									 -- x"7575547D", x"838E9A80", x"798387A0", x"91968382", x"967C919F", x"B8AD95A9", x"A7A8AF89", x"92257656",
									 -- x"24436DE0", x"C186CB7D", x"1D80756D", x"6D737DA2", x"B6877866", x"643683A8", x"C9B4BBBC", x"BFB6C1B1",
									 -- x"62263D93", x"52625A97", x"808A6675", x"85745783", x"7C7F7F6C", x"72988880", x"9385A3AE", x"A8B3A8A4",
									 -- x"B7A7B8B2", x"C79A604E", x"5F615A55", x"5756545B", x"52585C57", x"52515354", x"53535454", x"524F4F52",
									 -- x"4D4E4E4E", x"4C4A4847", x"44434240", x"3F3F3F3F", x"3F3C3A39", x"38373739", x"37353331", x"31313131",
									 -- x"2F2E2D2D", x"2C2C2D2D", x"2B2B2B2A", x"28272727", x"29282727", x"28292827", x"27282828", x"292B2B29",
									 -- x"2D2C2A2A", x"2B2C2D2D", x"2A2C2D2B", x"2B2E2E2C", x"2C2C2C2A", x"28292929", x"27262627", x"27272728",
									 -- x"27252424", x"24222021", x"23242626", x"25232120", x"24242324", x"24252627", x"27262729", x"2A29282A",
									 -- x"2C2C2B2B", x"2B2C2D2E", x"312F2D2B", x"2B2C2E2F", x"2A29302D", x"2C2F292D", x"2D353027", x"2127465B",
									 -- x"8BA3966C", x"87ABB7B4", x"B0AAAEA9", x"ADADADB5", x"A3A9A3A0", x"9CA0A9AC", x"AAACAFA8", x"A8ABA49D",
									 -- x"ECEBEBEA", x"EAEAEAEB", x"ECECEDEE", x"EEEEEDEC", x"EAEAEAE8", x"E7E7E7E7", x"E8E7E7E8", x"E8E8EAEC",
									 -- x"EAEBEBEA", x"EAEAEAEB", x"ECEBEBEB", x"EBEAE9E9", x"EAE9EBED", x"EEEDEDED", x"EFEFEFF0", x"EFEEEEEE",
									 -- x"ECECEDED", x"EDEDEDED", x"EDEEEFEF", x"F0F0EFEF", x"F0F0EFEF", x"EFEFEFEF", x"EFF1F2F1", x"EFEEEEF0",
									 -- x"F0F0EFED", x"ECECEAE7", x"E6E2DEDB", x"D5CECBCA", x"CDCDCDCD", x"CBC9C7C5", x"C2C2C1C3", x"C6C8C7C6",
									 -- x"C3C2C1C2", x"C2BEBBB9", x"BABCBFC2", x"C4C6C6C5", x"C7C6C7CA", x"CAC8C9CD", x"CDC8C3C0", x"BEBDBBB9",
									 -- x"BBBEBFBE", x"BEC0C1C0", x"BDB9B8BC", x"BBB8B9BD", x"BBBAB6B2", x"B0B0AFAF", x"AFADADAF", x"ACA5A2A3",
									 -- x"A6A6AAB0", x"B0ADB0B6", x"B3B4B4B4", x"B2AFADAC", x"A3ACB2AD", x"A7ABA99F", x"958E8D8A", x"88867F80",
									 -- x"77707E70", x"6B6D7493", x"7D5E6051", x"505B505E", x"5E564D61", x"545E5058", x"738F815C", x"5D4A232D",
									 -- x"5868649B", x"79577477", x"61336893", x"81723D69", x"876D635D", x"5B525844", x"2313565A", x"48565E7D",
									 -- x"4F2E3830", x"333F3B2E", x"40341E2B", x"4B798868", x"5F938564", x"9F9B967A", x"50679583", x"6E5B6969",
									 -- x"886F809B", x"7E48758E", x"847B8770", x"7280B396", x"A180918C", x"A9A5A197", x"AF8C9FB8", x"3B57C433",
									 -- x"71ABC690", x"7A98A8A7", x"353E7A56", x"70829168", x"4A3A0321", x"49333E4F", x"717A69B2", x"AD7FA0B0",
									 -- x"A45C2B48", x"3D717885", x"74537972", x"83777C7C", x"655A7595", x"6C829445", x"5C6BA079", x"8498919A",
									 -- x"A1A295A4", x"9FC0CA95", x"604B5462", x"58575D54", x"5E565256", x"59585759", x"52575954", x"4F52524D",
									 -- x"4C4D4E4E", x"4D4A4948", x"44454545", x"4443403E", x"403E3C3C", x"3B39383A", x"3A383635", x"34343434",
									 -- x"34333230", x"302F3030", x"2C2C2D2C", x"2A292929", x"29282828", x"28282827", x"2A2B2B2A", x"2B2C2C2A",
									 -- x"2C2B2A2B", x"2C2D2D2D", x"2D2F2F2D", x"2D2E2D2B", x"2E2E2D2B", x"29292929", x"2B2A2A29", x"28272727",
									 -- x"27252424", x"24222122", x"25252626", x"25232221", x"27272626", x"27272829", x"29292A2C", x"2C2B2B2C",
									 -- x"2D2E2F30", x"302F2E2E", x"26282B2E", x"302F2E2D", x"2A2A342D", x"292D2A34", x"292E2B4D", x"5B869096",
									 -- x"92A2B1AE", x"BAB5AAAC", x"B1B5A6AC", x"AFB3AABB", x"A197A3AC", x"AAA2A190", x"A5A19BAA", x"AF997B5B",
									 -- x"E3E4E4E5", x"E5E5E5E4", x"E9EAEBEC", x"EBEAE8E7", x"E7E7E7E6", x"E5E4E4E5", x"E4E4E5E7", x"E7E7E9EB",
									 -- x"EAEBEBEB", x"EAEAEBEB", x"ECECEBEB", x"ECECEBE9", x"EAE9EAED", x"EEEEEEF0", x"F1EFEEEE", x"F0F1F0EE",
									 -- x"EFEFEFEF", x"F0F0EFEF", x"EEEDEDEE", x"EEEFF0F1", x"F0F0F0F0", x"F0EFEEEE", x"F0F1F3F2", x"EFEDEEEF",
									 -- x"EFF0EEEC", x"EBECEBE9", x"EAEBECEB", x"E6DFDBDA", x"DAD9D9D9", x"DADADBDC", x"D3CFCCCC", x"CDCECDCC",
									 -- x"C8CACAC6", x"C5C6C2BB", x"BCBCBDC0", x"C2C4C5C6", x"C5C4C6CA", x"CBC9C9CD", x"CBCAC8C5", x"C3C3C3C4",
									 -- x"C3C3C2C0", x"BFC0C1C1", x"C1BFC2C7", x"C7C3C4C9", x"C7C5C1BC", x"BBBDBDBC", x"BEBDBBB9", x"B8B6B2AE",
									 -- x"B4B2B4BB", x"BDB9BABD", x"BDBEBFBE", x"BBB8B5B3", x"AFB2B6B5", x"B2B4B3AD", x"A0979490", x"90908886",
									 -- x"79797775", x"667C8B6D", x"65637973", x"66786F6C", x"5C60585B", x"665B6561", x"616B6161", x"54401C25",
									 -- x"5A5D8C7C", x"67757278", x"754F367C", x"75754A50", x"656E6C86", x"6A595C46", x"221F496C", x"49545963",
									 -- x"7F824D2D", x"48363712", x"2A3B2633", x"36235868", x"59686B7C", x"7A84868A", x"74535A70", x"7F8D9760",
									 -- x"7E809E86", x"838D9A86", x"9B8064AC", x"9D9BAAA8", x"9FA2A98B", x"93572B5F", x"7770B27E", x"68E08985",
									 -- x"C4B19B7E", x"5996BFA3", x"8D3C4E5C", x"5C3D3D37", x"576481DF", x"BEA691A5", x"8B818477", x"9E70904A",
									 -- x"66552F29", x"69485637", x"4569947C", x"777AA28C", x"6F807176", x"5A4A8186", x"6C57A492", x"A99EA997",
									 -- x"A8A19BA7", x"B9A7B5C1", x"C98B5550", x"5D5D5A5F", x"545C5E59", x"585B5A55", x"5F555354", x"5251514D",
									 -- x"4D4E4E4E", x"4D4B4B4A", x"47464747", x"47454240", x"41404042", x"413E3C3C", x"3B3A3938", x"38373635",
									 -- x"37363433", x"32323232", x"2D2D2E2D", x"2C2B2B2B", x"2C2B2B2A", x"2A2A2A29", x"2B2C2C2B", x"2C2D2D2B",
									 -- x"2B2A2A2A", x"2B2C2D2D", x"2F303130", x"2F2E2C2A", x"2E2D2D2C", x"2B2A2B2B", x"2E2E2D2B", x"2A292827",
									 -- x"28262626", x"26242426", x"25252526", x"27282829", x"29292929", x"292A2B2B", x"2C2C2C2E", x"2F2E2E2F",
									 -- x"2E2F3030", x"30302F2E", x"30302F2F", x"2F2E2E2E", x"362E302F", x"34362923", x"29346985", x"7F8F8F93",
									 -- x"9B929495", x"817A829C", x"A0AEB7AE", x"9BA2ACAF", x"ABA6A3A9", x"AEBABFC8", x"AC939D69", x"6A9B828C",
									 -- x"E0E1E2E3", x"E4E4E3E3", x"E4E5E6E7", x"E6E5E4E4", x"E4E4E5E4", x"E3E2E2E2", x"E1E1E2E4", x"E5E4E5E8",
									 -- x"EAEAEBEA", x"EAEAEBEC", x"EBEBEAEB", x"EBECECEB", x"EBEBECED", x"EDEBECED", x"EEEFEFEF", x"F1F2F0ED",
									 -- x"EFF0F0F0", x"F0F0F0F0", x"EEEDEDEC", x"EDEEF0F1", x"EDEEEFF0", x"F0F0EFEE", x"F1F2F3F2", x"F0EFEFF0",
									 -- x"EEEEEEEC", x"EBEDEDEC", x"ECEDEEED", x"EAE7E6E5", x"E4E4E4E4", x"E4E6E7E8", x"DEDAD7D7", x"D8D9D9D9",
									 -- x"D2D4D0C8", x"C6C9C6BD", x"BBBABABD", x"BFC1C3C4", x"C3C3C5C7", x"C8C8C7C8", x"C7C9CAC8", x"C5C4C5C7",
									 -- x"C7C7C8C7", x"C6C6C6C6", x"CACBCFD3", x"D3D0D2D5", x"D4D2CDC9", x"CCD2D5D3", x"D3CFC9C4", x"C2C1BEBA",
									 -- x"C4C2C3C8", x"CAC8C7C7", x"C5C7C9C7", x"C4BFBCBB", x"BEBBBCBC", x"B9B8B6B2", x"AAA39F9A", x"9B9D938E",
									 -- x"8D79756F", x"75876D75", x"73716686", x"737F7463", x"6865684E", x"77688147", x"4D605D52", x"3D1F274D",
									 -- x"65646E6E", x"676B6384", x"73761B5A", x"8C756234", x"68736B6A", x"572B745C", x"43392B5D", x"58544459",
									 -- x"39574833", x"393C2E27", x"1A2C1B13", x"2A302037", x"59455E72", x"6A6E5774", x"8C7AA178", x"7368875F",
									 -- x"64677B6E", x"6C716B89", x"859E738B", x"9591A59F", x"B1A57E6D", x"7B686196", x"8D8F6B43", x"5B8B7261",
									 -- x"9C889FA1", x"A095A9A3", x"AB77363A", x"4586B46C", x"CBB6ADB6", x"9AAA7F82", x"8A414542", x"41653453",
									 -- x"44725929", x"332F385C", x"69705177", x"797D717C", x"6F82A282", x"79797EA6", x"9E5E6082", x"AEAAA1AA",
									 -- x"B5B3AEB7", x"ABA595A9", x"ACCAB375", x"5452514F", x"595D5B53", x"51565B5B", x"5252595A", x"5152554F",
									 -- x"4F4F4E4E", x"4D4D4C4B", x"4C4A4847", x"47474645", x"41414244", x"43403E3D", x"3D3C3B3A", x"3A393736",
									 -- x"37363534", x"34343434", x"2F2F2F2F", x"2E2D2D2E", x"2D2C2C2C", x"2B2B2A2A", x"2B2C2C2C", x"2C2D2C2A",
									 -- x"2B2A2A2B", x"2C2D2D2D", x"2F303132", x"31302E2D", x"2D2D2E2F", x"2E2D2D2F", x"2E2F2F2D", x"2C2D2C2B",
									 -- x"2C2A2A2B", x"2A28292C", x"2B2A2A2A", x"2B2C2D2D", x"2B2B2B2B", x"2B2C2D2E", x"2F2E2F31", x"312F2F30",
									 -- x"302F2E2E", x"2E2F2F30", x"302F2E2D", x"2E303334", x"2C302E23", x"191E3448", x"739DA4A0", x"958E9AA0",
									 -- x"918A93A7", x"A7B6AFA5", x"9E95A5AC", x"B6A1A1B3", x"ADB8B4AF", x"939C7D65", x"81878180", x"8C9FA9A0",
									 -- x"E0E1E1E2", x"E3E4E4E4", x"E2E3E2E1", x"E0E0E1E2", x"E2E3E4E4", x"E3E2E1E1", x"E0E0E1E2", x"E2E2E3E5",
									 -- x"E8E9E9EA", x"EAEAECED", x"EAEAEAE9", x"E9EAEAEB", x"EBEBECED", x"ECEAEAEC", x"ECEEEFEE", x"EDEEEFED",
									 -- x"EFEFEFEF", x"EFEFEFEF", x"EEEEEDED", x"EDEDEEEE", x"ECEDEDEE", x"EEEFEFEF", x"F1F2F3F2", x"F1F0F0F1",
									 -- x"EEEFEEEC", x"ECEEEEEE", x"EDEDEDED", x"ECECEBEB", x"ECEDEEEF", x"EFEEEEED", x"E7E4E1E2", x"E2E0E0E1",
									 -- x"DBDAD5CE", x"CBCCC7C0", x"BAB8B8BA", x"BCBCBBBC", x"BFC1C2C3", x"C4C5C5C3", x"C3C5C7C7", x"C4C3C4C6",
									 -- x"C7C8C9CA", x"CAC9CACB", x"CDD1D6D8", x"D8D8DADD", x"D6D7D7DA", x"E3EFF3F1", x"E4DDD6D1", x"CCC7C5C6",
									 -- x"D0D1D3D5", x"D6D5D4D3", x"D1D3D5D5", x"D1CCC9C8", x"CCC9C8C5", x"BFBDBAB5", x"AFACABA3", x"A4A79C95",
									 -- x"8C82807D", x"7A7F6E57", x"6E755B63", x"857A6D68", x"5B63627C", x"6B676555", x"7087355C", x"56575144",
									 -- x"60867977", x"455A7267", x"7B6A4132", x"5C7A4F70", x"95705257", x"48679085", x"53685C3F", x"2C4A2C05",
									 -- x"3E3A4A23", x"1512162E", x"22191C43", x"55645D60", x"5C586473", x"7A566B95", x"7F82838A", x"57091E48",
									 -- x"4338505A", x"585B6360", x"4B928984", x"A38B9787", x"8D7D8F88", x"947B5974", x"6A3D1843", x"12052866",
									 -- x"6E818093", x"C39498B4", x"99813738", x"2C94885B", x"4F404877", x"8BA17D87", x"60642C6E", x"61706B4F",
									 -- x"67B6733A", x"1D352047", x"37896C6E", x"9C8C8393", x"8D8A946F", x"9B7B84A1", x"9587D592", x"9296ACA8",
									 -- x"9C75B9A3", x"A3A2899D", x"8E8CB4C8", x"A498AFB5", x"5E4F5A7E", x"8D775C53", x"53545D5D", x"53565A53",
									 -- x"53525151", x"51504E4C", x"504D4A49", x"494A4948", x"44434344", x"43413F40", x"41403E3D", x"3C3B3A39",
									 -- x"39393837", x"36363535", x"33333231", x"302F3030", x"2D2E2D2D", x"2C2B2B2B", x"2C2D2D2D", x"2D2E2D2B",
									 -- x"2D2D2C2D", x"2E2F2F2F", x"30313233", x"33323130", x"302F3032", x"322F2F30", x"2F30302E", x"2E302F2E",
									 -- x"302F2E2F", x"2D2C2D30", x"302F2D2D", x"2D2D2C2B", x"2C2C2C2C", x"2D2E2F30", x"31303132", x"32303031",
									 -- x"31302F2F", x"2F303132", x"35343331", x"2E2A2624", x"23333F5A", x"6F7A8D8E", x"6E9691A2", x"90999FAF",
									 -- x"A79496A5", x"B1BBBEC4", x"ADB4B49A", x"8C6D5A7E", x"91544E7D", x"7649314E", x"7A809DBC", x"AA7B6F82",
									 -- x"DFDFDFDF", x"E0E1E3E4", x"E3E2E0DD", x"DCDCDEE1", x"E1E2E4E4", x"E4E2E1E1", x"E2E1E1E2", x"E1E1E2E5",
									 -- x"E7E7E8E9", x"E9EAECED", x"ECECECEA", x"E9E9EAEB", x"EAEAEDEF", x"EFEDECEE", x"ECEFF0EC", x"E9EBEEF0",
									 -- x"F1F0F0EF", x"EFEFEFEF", x"EEEEEEED", x"EDECECEC", x"EDEDECEC", x"ECEDEEEF", x"F1F1F2F2", x"F1F0F0F0",
									 -- x"EFF0F0EE", x"EDEEEFEE", x"F0F0F0F0", x"F1F1F0EE", x"EDEFF3F6", x"F7F6F5F3", x"EEEBE8E7", x"E4DFDCDC",
									 -- x"DDDAD6D3", x"D1CCC6C1", x"BAB8B7B9", x"B9B6B4B4", x"B8BCBDBD", x"BFC2C2BE", x"BEC1C4C6", x"C6C6C8C9",
									 -- x"CACAC9C8", x"C7C7C8C9", x"CBD0D5D6", x"D6D9DDDF", x"E5E6E8EB", x"F3FBF9F3", x"E9E1DDDD", x"D8CECCD2",
									 -- x"D4D8DBDB", x"DBDBDBDA", x"DCDFE2E1", x"DED9D6D5", x"D3D3D3CE", x"C8C7C5BE", x"B9BBBCB4", x"B2B6ABA2",
									 -- x"9E888776", x"7A736672", x"7783755B", x"48686B65", x"4676716F", x"656F6C85", x"72676150", x"4163625C",
									 -- x"6C7A7469", x"69766E6E", x"646F5E32", x"59456278", x"676A5D7A", x"4B669592", x"297F894D", x"240B0C29",
									 -- x"212E2E5B", x"503D2929", x"65709199", x"9EA58898", x"703C4563", x"6F59618A", x"7D7D7172", x"7F5B1C26",
									 -- x"254C593D", x"4C445F4A", x"3D8D8683", x"7E7A868C", x"8BAA8A66", x"A390823D", x"1A010202", x"0935638C",
									 -- x"94869EA7", x"ADABC1B5", x"945E283F", x"72502322", x"1B230D17", x"815A4957", x"8285926C", x"43899C6B",
									 -- x"5B919845", x"28506A48", x"30578338", x"53A5846E", x"77806C76", x"8B7F9194", x"76795A97", x"8885A49B",
									 -- x"A8A4C29F", x"938DADAE", x"B19586A1", x"BFBAB1BE", x"96A9B9C0", x"C9CEBFA8", x"79584F5B", x"5C585A58",
									 -- x"5A585757", x"5756524F", x"504F4D4D", x"4E4D4B48", x"49474545", x"44434344", x"4644413F", x"3E3D3D3C",
									 -- x"3D3D3C3A", x"39373635", x"35353432", x"31303132", x"30303030", x"2E2E2E2E", x"2D2E2F2E", x"2F302F2C",
									 -- x"2F2F2F2F", x"30313130", x"33323233", x"33323232", x"33333335", x"33302F30", x"3031312F", x"2F31312F",
									 -- x"32313130", x"2F2D2E31", x"2C2C2C2D", x"2E2E2C2B", x"2C2C2C2C", x"2D2F3031", x"33323233", x"33313031",
									 -- x"30313233", x"34333332", x"312C2626", x"2E3F515C", x"759199A5", x"9B8EA1A4", x"702E9C9D", x"A6909697",
									 -- x"969BA195", x"A1ABB2B7", x"AB9A837E", x"81AC959A", x"B5BAB28B", x"A9A7BCE6", x"C4A7A888", x"8B9E7367",
									 -- x"E0E1E1E1", x"E1E1E2E3", x"E1E0DEDE", x"DEDEDFDF", x"E1E0E2E5", x"E5E3E1E2", x"E3E2E1E2", x"E3E5E5E5",
									 -- x"E8E8E8E9", x"E9E9EAEA", x"EDEBEAEA", x"EBEBEBEA", x"EAEAEBEC", x"EDEDEDED", x"EEEFEFEF", x"EDEBEAE9",
									 -- x"EEEEEFEF", x"EFF0F1F2", x"EFEFEEED", x"EDEDEDED", x"EDECECEE", x"EEEEEEF0", x"F2F2F2F1", x"F0F0F0F1",
									 -- x"F0EFEDEC", x"EDEFF0F1", x"F0F0F0F0", x"F0F0F0F0", x"F1F2F3F5", x"F7F8F8F8", x"F5F0ECE9", x"E5E0DDDD",
									 -- x"D9D9D7D4", x"D1CEC8C2", x"BDB6B3B4", x"B4B4B3B0", x"B6B5B6B7", x"B6B5B8BD", x"C1BFBFC1", x"C3C2C1C2",
									 -- x"C5C3C4C7", x"C7C4C5CA", x"CACDD1D4", x"D6D9DDE0", x"E4E8EAED", x"F3F7F3EB", x"E6DCD8D8", x"D3CECFD1",
									 -- x"D3D7DBDD", x"DFDFE0DF", x"DFE3E5E3", x"E0DFDDDB", x"D8D7D6D1", x"CAC9C9C5", x"C4C5C7C6", x"C3C0B7A9",
									 -- x"9D948B7D", x"73587485", x"7573767E", x"717A616F", x"6B8D786B", x"69647559", x"65594A5D", x"56696365",
									 -- x"6B75787B", x"64767173", x"7D757D4A", x"4B8A7869", x"706B566F", x"2D596C57", x"398C7390", x"8A6E3F1F",
									 -- x"1A102F89", x"7E7754A7", x"A1A2897C", x"787C7480", x"92B2712B", x"40464030", x"2D374B35", x"437F713B",
									 -- x"3D2B4843", x"414F585D", x"495D6E66", x"848B59A4", x"9A75807E", x"772D0300", x"1B24282E", x"434E6B8C",
									 -- x"8C9FD2A7", x"988C9DAB", x"AB921C1B", x"7DB09B60", x"455F2E35", x"5B57B8AE", x"9DA6A76D", x"5D6C9EA5",
									 -- x"58576C72", x"401C4E54", x"6867354A", x"437C7069", x"77698B7F", x"A1B5AF68", x"89859272", x"7A675A92",
									 -- x"AEB57F90", x"99938A8F", x"9DA9988B", x"A09FADB7", x"B6A895A4", x"A4ADB2C6", x"CAA96A48", x"57665E5B",
									 -- x"5B63585A", x"5C5C5255", x"53525053", x"5250534F", x"504B4747", x"4A4B4946", x"45474644", x"42413F3C",
									 -- x"3D3C3B3A", x"3A3A3938", x"36373533", x"33353330", x"3034322C", x"33342D35", x"342C2C31", x"312F3031",
									 -- x"372C3138", x"2D2C3437", x"333C3932", x"3D343537", x"34323633", x"32332F31", x"31363031", x"30322E34",
									 -- x"2A2D3131", x"302F3032", x"332B2A2E", x"302F2F2E", x"2C2E2D32", x"302A3835", x"35353335", x"36343234",
									 -- x"372E303D", x"35313233", x"343D6867", x"A59FB4B7", x"9CAC9E9E", x"9580AEAA", x"9E225B9D", x"998C7192",
									 -- x"989AA1A5", x"A9AAAF9F", x"8A8BA6BE", x"CDC1BEA2", x"939A8C68", x"66A19389", x"84687879", x"78576A49",
									 -- x"DDDEDFDF", x"DFDFDFDF", x"E0DFDFDE", x"DFE0E0E0", x"E2E1E2E4", x"E4E2E1E2", x"E3E3E3E4", x"E4E5E5E6",
									 -- x"EBEAEAEA", x"EAEBEBEC", x"ECEBEAEA", x"EBECECEC", x"EDEDEDEE", x"EEEEEEEE", x"EFEFEFEE", x"EDEBEAEA",
									 -- x"EEEFF0F1", x"F1F0F1F1", x"F0F0EEED", x"EDEDEDEE", x"F0EEEEEF", x"EFEEEFF1", x"F3F3F3F3", x"F2F2F2F3",
									 -- x"EFEEEEEF", x"EFEFEFEE", x"F0EFEFEF", x"EFEFF0F0", x"F1F1F2F4", x"F6F7F8F7", x"F7F3F0EE", x"EAE4DFDD",
									 -- x"DBD9D6D3", x"D2D0CAC5", x"BEB7B4B4", x"B1B0B2B0", x"B0AFB0B1", x"B2B3B7BC", x"BEBBBABB", x"BDBDBEC0",
									 -- x"BFBEBFC1", x"C0BDBFC4", x"C7C8CACE", x"D4D8DBDC", x"E2E4E6E8", x"EDF0ECE5", x"DFD1CBCF", x"D0CFCFCE",
									 -- x"D4DBDFDD", x"DDDFDFDB", x"DFDFDFE0", x"E2E2DCD5", x"D6D5D6D3", x"CDCDCECA", x"CAC9CBCC", x"CBC9BEAF",
									 -- x"A49C997A", x"6D69776B", x"79746985", x"71696476", x"747A8472", x"5B846350", x"57635567", x"917E5961",
									 -- x"88706E93", x"7E7C9079", x"836C4C6D", x"58787980", x"6E676080", x"38557159", x"36636971", x"6B71733A",
									 -- x"281D3F68", x"794E7E93", x"69769095", x"7C6E6F6B", x"98614384", x"5C3B5B28", x"021F2E39", x"3F63272C",
									 -- x"9D260302", x"343C2C3A", x"5762737F", x"9E9A8C8B", x"658A8487", x"AD28415E", x"7CAE835F", x"546477BA",
									 -- x"8C89A68B", x"AF979EA9", x"B2803017", x"5ECA4B4F", x"8C385250", x"1698B297", x"94909FA9", x"8C91AF8F",
									 -- x"887F6F7C", x"97381033", x"4E6F6F8D", x"6871727E", x"8C7B868D", x"96968773", x"86878F97", x"8F99BBA8",
									 -- x"B9AFB2BB", x"A5A3677D", x"8A8A9193", x"9891C3C4", x"B1B79A8C", x"A7A4A9B0", x"BBA9BB8C", x"795A4B58",
									 -- x"5E606065", x"5F5B5D5D", x"5B5C5B5C", x"58535453", x"504E4B4A", x"4B4B4A49", x"47484745", x"44454442",
									 -- x"3D3E4041", x"413F3B39", x"3D3A393A", x"3A383839", x"37393C38", x"39352E35", x"31353630", x"2F37382D",
									 -- x"2E353234", x"343A3331", x"343A343C", x"323A3737", x"39343635", x"36373233", x"2E363332", x"3739302C",
									 -- x"31303030", x"30302D2B", x"2B31342F", x"2C2D2E2D", x"2F33322A", x"32342823", x"212B2A2D", x"2D384036",
									 -- x"323E3426", x"272A322A", x"2687CB85", x"65A2A09C", x"A09C9FA3", x"B7A58F8B", x"815A218B", x"9DA46579",
									 -- x"9A7891B5", x"BFA1AAC2", x"AAC2B395", x"93908F52", x"4A486871", x"71793920", x"4B604C4D", x"54575F57",
									 -- x"DCDDDEDE", x"DEDEDFDF", x"DFDFDEDE", x"DEDEDEDD", x"E1E0E0E2", x"E2E2E2E4", x"E5E6E7E7", x"E7E6E7E8",
									 -- x"ECEBEAEA", x"EAEAEBEC", x"ECEBEBEC", x"EDEEEEEE", x"F1F0F0F0", x"F0EFEFEF", x"EFEFEFEE", x"ECEBEBEC",
									 -- x"EFF0F1F2", x"F2F1F0F0", x"F0EFEEED", x"EDEEF0F0", x"F2F0EFEF", x"EFEEEFF1", x"F4F4F4F3", x"F1F0F0F1",
									 -- x"F1F1F0EF", x"EFEFEEEE", x"EFEFEFEE", x"EEEFEFEF", x"F1F1F2F3", x"F6F7F8F8", x"F6F5F4F4", x"F0E9E3E0",
									 -- x"DEDBD6D3", x"D3D1CBC5", x"BFB9B5B3", x"AEADB0B0", x"AFADABAC", x"ADAFB2B6", x"B9B6B5B6", x"B8B8BABB",
									 -- x"BAB9BABC", x"BAB8BBBF", x"C2C1C2C8", x"CFD5D8D7", x"DFE0E1E2", x"E7EAE7E2", x"DCD0CCD1", x"D3D3D3D1",
									 -- x"D3DBDED9", x"D9DFE1DD", x"E1E0E0E1", x"E3E2DBD3", x"D4D3D6D5", x"D2D2D3D0", x"CDCACBCD", x"CECDC3B3",
									 -- x"B4AD8D69", x"7576715B", x"4A697C58", x"6B73697A", x"6B8B7F5E", x"6A6C6860", x"81896C7E", x"7D6E4622",
									 -- x"2C58636B", x"7C6A6B71", x"6C576B8F", x"416A9974", x"4D618A77", x"1A6F8360", x"66756658", x"737A7064",
									 -- x"3A5B4E55", x"6E4E7D8F", x"77747871", x"62628562", x"4D6B8079", x"8483A079", x"361A2314", x"1C210253",
									 -- x"7EB58D22", x"00000814", x"0F101C37", x"4E867358", x"777979B7", x"751BA08D", x"B99D795D", x"5C8A72C2",
									 -- x"9DADC198", x"936BB1A9", x"AE5E411E", x"559A3D64", x"ABA59774", x"0D89696F", x"919C93B6", x"968F866A",
									 -- x"73607F76", x"7F971C53", x"96805D59", x"735D706C", x"8C829C89", x"847B856C", x"9287708F", x"A3C5E0A1",
									 -- x"9A89C2B6", x"9E9F8F65", x"636988AC", x"968190A2", x"A8A8BD9F", x"7C99A9B9", x"B9C28E6B", x"B9B79584",
									 -- x"725A5769", x"626F6761", x"625E5B5A", x"5A585554", x"52535351", x"4E4C4D4E", x"4C4C4B48", x"47474645",
									 -- x"44434241", x"42424242", x"423E3D40", x"3F3B3B41", x"40373635", x"383B383D", x"37363737", x"35383834",
									 -- x"41353C38", x"372D3A3C", x"38373634", x"3A3C3C3A", x"3A363836", x"36363336", x"39303536", x"2C2C3736",
									 -- x"3131312F", x"2F303437", x"2F302F2F", x"32312E2F", x"33363037", x"2C32477E", x"88767969", x"3829273B",
									 -- x"35214A6C", x"91A1A49B", x"7D3D7CAF", x"586A9A5A", x"7F938398", x"7F59334D", x"75783F0D", x"93A4824B",
									 -- x"7F724166", x"79965944", x"9FC9BC8A", x"515B8184", x"8D909299", x"A98D5A62", x"6D8C808B", x"91875E78",
									 -- x"E2E2E3E3", x"E3E4E5E7", x"E3E2E1E1", x"E0DFDEDD", x"E0E0E1E3", x"E4E5E6E7", x"E8EAECEC", x"EAE9EAEC",
									 -- x"EDEDECEC", x"ECECEDED", x"EEEEEEEF", x"F0F1F1F1", x"F3F3F3F2", x"F2F2F2F1", x"F0EFEFED", x"ECECEDEE",
									 -- x"F0F1F2F2", x"F1F1F0F0", x"F1F0EEEE", x"EFF0F2F4", x"F2F0EFEF", x"EFEEEFF1", x"F3F3F4F4", x"F3F3F3F4",
									 -- x"F8F6F3F0", x"EEEEEFF1", x"F0EFEFEE", x"EEEEEEEE", x"F0EFF0F1", x"F3F5F6F6", x"F3F4F5F6", x"F4EEE8E4",
									 -- x"E2DFDAD7", x"D7D4CCC3", x"C2BAB6B4", x"AFAEAFAE", x"AEACA9A9", x"AAADAFB0", x"B2B1B1B4", x"B5B5B6B7",
									 -- x"B7B4B4B5", x"B6B6B8BA", x"BAB9BBC0", x"C7CDD0D0", x"D8D9DADC", x"E2E6E6E2", x"D6D0D1D4", x"D2CFD0CF",
									 -- x"D5D8D8D4", x"D4DADFE1", x"DDE0E1DF", x"DAD6D2D1", x"CECED2D4", x"D2D3D4D1", x"D1CECFD1", x"D2D2CBBF",
									 -- x"BDBA8680", x"83779264", x"75997D6A", x"6B767D71", x"9B6E7C8C", x"80884965", x"7C6E7B74", x"5B530A33",
									 -- x"343A644D", x"5C634D63", x"4C4F5253", x"18477858", x"70636B4F", x"1E616067", x"74697687", x"6F7D867F",
									 -- x"41708A63", x"374B5923", x"364E4B38", x"4F4A552C", x"66987070", x"6E727C61", x"6F20090E", x"1E064383",
									 -- x"92959F55", x"1E3B0F06", x"00040000", x"0D294753", x"48708599", x"3A4887A6", x"95B5988A", x"697B8FB2",
									 -- x"95B58D8A", x"B79666AC", x"8F710123", x"A782586E", x"6A77739A", x"702A4624", x"4373A59B", x"A9A57055",
									 -- x"8CAF807C", x"59837CB6", x"BCB8A67A", x"507C7E6D", x"75876D8A", x"8A8D637E", x"AD917F82", x"8F989C93",
									 -- x"8F919588", x"9C7A608D", x"7F947F87", x"9F9F849C", x"B48394CA", x"BA925F5C", x"6970915C", x"6391A7A2",
									 -- x"D7D2A07A", x"6460696B", x"66636460", x"5E5E5B5A", x"58595957", x"54525354", x"5252504E", x"4D4C4B4B",
									 -- x"4E4C4947", x"46474747", x"46434244", x"423F4146", x"413C3F3E", x"3C3D3937", x"4039393D", x"3A36373A",
									 -- x"2D393336", x"3D342531", x"474E5243", x"4C392A27", x"2A2C3536", x"36363439", x"3D373839", x"39353532",
									 -- x"34353635", x"33302E2E", x"34332F30", x"36363334", x"30363524", x"407AAF9B", x"8C809FAB", x"96905F45",
									 -- x"45789DB7", x"A39496B5", x"C1A75031", x"8935409F", x"167B7A2E", x"7697AA8F", x"A297AA35", x"218072AB",
									 -- x"7E80818A", x"A4A6BC54", x"306C7A57", x"53A6ADC1", x"C5D4ACA6", x"BA9A97A2", x"9796A5A5", x"8F9F9F8F",
									 -- x"EAEAEAEA", x"EAEBECED", x"E9E9E8E8", x"E7E7E5E4", x"E3E4E6E7", x"E9EAEBEA", x"ECEEF0F0", x"EEEDEEEF",
									 -- x"EFF0F0F1", x"F1F1F0F0", x"F1F2F2F3", x"F3F3F3F4", x"F5F4F4F4", x"F3F4F4F4", x"F2F2F1F0", x"EFEFF0F1",
									 -- x"F4F4F4F4", x"F3F2F2F3", x"F3F2F1F0", x"F0F2F4F5", x"F3F1F1F2", x"F2F2F3F5", x"F3F5F7F9", x"FAFBFDFE",
									 -- x"FDFCF8F4", x"F1EFF0F1", x"F0F0EFEE", x"EEEDEDED", x"EDEDEDEE", x"F0F2F3F3", x"F2F4F5F6", x"F5F1EDE9",
									 -- x"E6E4E0DE", x"DEDAD0C7", x"C4BCB7B6", x"B2B1AFAC", x"A9A7A6A6", x"A9ACADAD", x"ABAAABAD", x"AFB1B3B7",
									 -- x"B2AEACAE", x"B2B4B4B4", x"B2B3B6BA", x"BFC3C7C9", x"CDCED1D5", x"DDE2E3E2", x"D5CFCFD2", x"D1D1D4D4",
									 -- x"D7D3D1D2", x"D3D3D8DE", x"D7D8D9D4", x"CDC7C7C9", x"C5C5CACF", x"CFD1D2D0", x"CFCDCFD1", x"D1D2D1CA",
									 -- x"D7A0795D", x"6C7E7371", x"8081636B", x"9161737B", x"6A80827D", x"746B6780", x"8B777F7A", x"8B752932",
									 -- x"787D5C4F", x"4A55825D", x"593C3A3F", x"246E4D63", x"7E906C3D", x"697C8476", x"6F847378", x"73807C7D",
									 -- x"5825848B", x"5F274A44", x"43132D19", x"1E41768A", x"86776664", x"67787662", x"48001B4A", x"4E3C2E2B",
									 -- x"46273F37", x"44906554", x"6344373A", x"1F0F0640", x"585D897F", x"616DA573", x"8FD18A93", x"929D8580",
									 -- x"63737481", x"73958A6E", x"71653561", x"857C6580", x"9E988F88", x"4C42101B", x"271852B9", x"B0A8C397",
									 -- x"A09B9378", x"7A52736B", x"BCA7B395", x"00384878", x"5F627570", x"8474796F", x"7F7A8F79", x"85918D9A",
									 -- x"97A18368", x"806CA594", x"A2B7A79C", x"8C93AC91", x"ABB29DA5", x"AEB73A6B", x"74A2E8DB", x"C8854B2B",
									 -- x"53B1DCD4", x"CCAE8C62", x"65606A68", x"60646465", x"5F605F5E", x"5C5B5A5A", x"59585757", x"56555454",
									 -- x"52535353", x"514D4845", x"4A4B4A47", x"45464748", x"42444A43", x"3C3F4041", x"403F403D", x"393B3E3C",
									 -- x"3F383D2E", x"27448DB8", x"D0CBBCAD", x"928C7675", x"675D5343", x"39393639", x"2F3F3A33", x"3C3B353E",
									 -- x"3D393434", x"37393937", x"31373935", x"34353534", x"2F2B1F35", x"4B5B4F63", x"9E9898A5", x"9CA6B5AE",
									 -- x"98977239", x"A19F90A1", x"90A3B74F", x"02101E5F", x"762E798F", x"A7B8B99E", x"B3ADA4CC", x"4F067FC3",
									 -- x"A193BCB4", x"A4A5B7CA", x"821150A9", x"B7A7A2CD", x"B3B6A09F", x"A594A48E", x"7691948B", x"94A2B3A1",
									 -- x"E8E9EAEA", x"EAEAEBEB", x"EBEBEAEB", x"EBECECEB", x"E9EBECEC", x"EDEEEEEC", x"EEEFF1F1", x"F0EFF0F1",
									 -- x"EFF0F1F2", x"F3F2F1F1", x"F3F4F5F5", x"F5F4F4F5", x"F5F5F4F4", x"F4F4F5F5", x"F4F4F4F3", x"F3F3F4F5",
									 -- x"F7F7F7F6", x"F5F5F6F7", x"F6F5F4F3", x"F2F3F4F5", x"F6F5F5F7", x"F8F8F8FA", x"FAFBFDFE", x"FEFEFFFF",
									 -- x"FEFEFDFA", x"F5F1EFEE", x"F0EFEEED", x"EDECECEC", x"EEEEEEEF", x"F1F2F2F2", x"F3F4F5F5", x"F4F2EFEB",
									 -- x"E9E7E5E4", x"E3E0D8D0", x"C7BEBAB8", x"B5B3B0AA", x"A7A6A4A3", x"A4A6A6A5", x"A6A4A3A4", x"A6A9AFB4",
									 -- x"ADAAA8AA", x"AEB0B0AE", x"AEB1B5B8", x"BBBEC2C5", x"C6C7CCD2", x"DAE0E1E1", x"D7CDC8CC", x"D1D9DDDC",
									 -- x"D2CBCACF", x"D2CFD2D9", x"D4D0CBC7", x"C4C1C0C1", x"BDBCC2CA", x"CCCFD1D0", x"CBCACDCF", x"CDCFD1D0",
									 -- x"CC814E62", x"6E6A8287", x"64737384", x"7C75758F", x"6989756F", x"7A777073", x"A6886175", x"59698639",
									 -- x"5A835741", x"3E55624A", x"5845600D", x"3B4F4361", x"6C704457", x"6D82776B", x"97788862", x"6F945A68",
									 -- x"7451626D", x"877C7968", x"6A887447", x"2D215B76", x"58474D4C", x"5F6A6588", x"2F050022", x"2F3A3D2D",
									 -- x"1B242700", x"3A958E96", x"859EAEAA", x"B6878D4F", x"2E253E68", x"918892A9", x"8C8F9C7A", x"B0AC86B1",
									 -- x"A492BB92", x"48625B7E", x"907B4865", x"AFBA946C", x"CBA2AB95", x"7E7D5E4D", x"59780946", x"ABC5BA87",
									 -- x"9A98947C", x"B8C6822D", x"AEAD844C", x"8EA38B58", x"5C466274", x"6B6B8A78", x"84787261", x"83807683",
									 -- x"9372719F", x"A0C0BA91", x"A27AAD8C", x"B07E808C", x"A0A5697E", x"A7B05F78", x"D4B3AAC5", x"CFD9BEA4",
									 -- x"4C52CCB2", x"C5C9D2BD", x"86656970", x"6C706C67", x"69686665", x"65656463", x"64625F5D", x"5B585758",
									 -- x"55555555", x"5553504D", x"4E4F4E4A", x"48494A48", x"47464741", x"41454141", x"3F3D3E3E", x"38343534",
									 -- x"2F2D3A62", x"99B79A68", x"5D48576A", x"7DAABFBE", x"BDB2A184", x"6E614C3F", x"42333541", x"30323739",
									 -- x"3B3C3D3B", x"37343333", x"392F3239", x"35303132", x"34619382", x"323F5295", x"9964675D", x"6C857487",
									 -- x"A994786D", x"809F996D", x"707095B8", x"674D4762", x"A6721B8D", x"7C69849E", x"646F7F48", x"B86A1F48",
									 -- x"A0AEACA2", x"ADA4AFB0", x"B8CF7BAD", x"B8AEB7AB", x"A39A9A94", x"9C9FA6AB", x"88A0B5A3", x"A5ACA09A",
									 -- x"DEE1E4E6", x"E7E7E7E7", x"E9E9E8E9", x"EAEBECEC", x"ECEDEDEC", x"EDEEEFED", x"EEEEEEEF", x"EFF0F0F1",
									 -- x"EFEFF0F1", x"F2F2F2F1", x"F3F4F5F5", x"F5F4F4F5", x"F5F5F4F4", x"F4F4F5F5", x"F4F4F4F4", x"F4F4F5F6",
									 -- x"F7F8F8F8", x"F7F7F7F7", x"F7F7F6F5", x"F4F5F6F6", x"FAF9FAFC", x"FDFDFDFE", x"FEFFFFFF", x"FFFDFDFC",
									 -- x"FDFEFEFA", x"F5F1EEED", x"EDEDECEC", x"EBEBEBEB", x"EEEEEFF0", x"F1F1F1F0", x"F0F2F3F2", x"F2F2EFEC",
									 -- x"EBE9E6E4", x"E4E3DED9", x"C9C1BDBB", x"B5B1AFAA", x"A8A7A4A0", x"9EA0A09F", x"A2A0A0A0", x"A1A2A6AA",
									 -- x"A7A7A6A7", x"A8A9AAA9", x"AAADB2B5", x"B7B9BCBF", x"C3C5CAD1", x"D7DBDCDC", x"D4C9C5C8", x"CED7DDDC",
									 -- x"D1C9C5C8", x"CBCBCDD1", x"CBC4BCB9", x"B9B8B7B6", x"B4B3B9C2", x"C6C9CCCB", x"CBCACCCD", x"C9C9CCCB",
									 -- x"C57B7F9F", x"7969807B", x"85615167", x"68746930", x"5F887E63", x"916A3F22", x"5470504B", x"3E55658F",
									 -- x"49705D87", x"7A775E58", x"5B0E002E", x"5356646D", x"8C514756", x"766F7A5C", x"76727581", x"84727366",
									 -- x"6B6A4F7D", x"71857B82", x"80728588", x"80673F46", x"4B174C24", x"454A4D5D", x"1900010D", x"25231F1B",
									 -- x"3A342654", x"7E7D948F", x"8A8F9CA2", x"9C8B9083", x"8B590966", x"7AA47E7C", x"8985868F", x"A3CBA8B4",
									 -- x"BEACBD74", x"064385D0", x"C5985C65", x"B8B5A694", x"6E71AB9C", x"AA9AA499", x"9B54092C", x"5B6789BC",
									 -- x"C58DC5B6", x"C396A0B8", x"6E5D7FB6", x"BEB5A9B0", x"714D4856", x"39697D41", x"55573B12", x"183D7589",
									 -- x"766F8BAD", x"9992B1B5", x"B998749D", x"7A3D3450", x"66725300", x"3768906F", x"87C69893", x"B7BFBCC5",
									 -- x"D3545BA8", x"BBC0A3C3", x"E3947B7B", x"6E6E7072", x"73727170", x"6F6F6F70", x"706C6764", x"605D5D5F",
									 -- x"5E5C5A58", x"58595959", x"5452504F", x"4D4B4A4A", x"4A494A49", x"4C463C43", x"3E424E59", x"5A5A5E60",
									 -- x"826E77A0", x"58555F79", x"5A608D9D", x"AFA58B72", x"313F5057", x"6C8EA2AB", x"A4807A8E", x"67625035",
									 -- x"2F33383C", x"3E3C3936", x"34373F35", x"24458EC1", x"A678B2AE", x"43013660", x"5854343B", x"68738065",
									 -- x"685E3369", x"5D436A7D", x"7B545131", x"67632C84", x"513F7F42", x"5C6067A1", x"90792242", x"8AA67A4D",
									 -- x"256E988F", x"A69A94A7", x"A0A5CDBE", x"9F78A4A6", x"888D9D9B", x"A28A6675", x"6090B7A8", x"B1AAA298",
									 -- x"D7DBE1E6", x"E9E9E9E8", x"E9E8E7E7", x"E8E9EAEA", x"EBECECEA", x"EAEDEFEE", x"EDEDECED", x"EEEFF0F0",
									 -- x"F0F0F1F1", x"F2F3F4F4", x"F1F3F4F5", x"F4F3F4F4", x"F6F5F4F3", x"F3F4F4F5", x"F2F3F3F3", x"F3F3F4F5",
									 -- x"F6F7F8F8", x"F8F7F6F6", x"F6F6F6F6", x"F6F7F8F8", x"FBFBFDFF", x"FFFFFFFF", x"FDFFFFFF", x"FFFFFFFF",
									 -- x"FEFEFCF8", x"F3EFEEEF", x"EBEBEBEB", x"EBEBEBEB", x"ECECECED", x"EEEEEDEC", x"ECEEEFEF", x"F0F1EFEC",
									 -- x"ECEAE6E2", x"E1E1E0DD", x"CAC3BFBC", x"B4AFAEAB", x"A5A5A29D", x"9C9EA0A0", x"A0A0A1A2", x"A09E9E9F",
									 -- x"A0A2A3A2", x"A1A1A2A3", x"A3A6AAAE", x"B1B3B5B7", x"C1C3C7CE", x"D4D6D6D5", x"D6D1D0D2", x"D2D7DDDE",
									 -- x"D9D0C6C1", x"C2C5C7C8", x"BDB6B0AC", x"AAA8A8AA", x"ACAAB0B9", x"BDC0C2C2", x"C3C0C1C1", x"BCBABBB9",
									 -- x"8F80756C", x"7C7D5D67", x"61484876", x"907A234E", x"65605285", x"5D4B4340", x"6642371B", x"114A666E",
									 -- x"6C99839B", x"64440004", x"0001506B", x"7CA3675D", x"5C51336F", x"7A757E75", x"6C6C677A", x"77646E6C",
									 -- x"6A795863", x"4F6E7373", x"7D8B7677", x"697B8F6E", x"66332754", x"49324F39", x"020B0C5F", x"968DA39A",
									 -- x"828F8479", x"81907F82", x"89939999", x"94918994", x"80816D01", x"003A6279", x"8298A6AD", x"B3A7B394",
									 -- x"8F83C534", x"2383CEB1", x"614B31AD", x"B1A0BAC8", x"80A8A49C", x"98A9A09F", x"B2964577", x"14092263",
									 -- x"8599BBCA", x"9D5066AB", x"7F35D5A7", x"A69F9AA4", x"BDAF744D", x"5B432F2D", x"321B588B", x"39002C4C",
									 -- x"59607682", x"8E94A1AA", x"D3B7AFBB", x"D3CDA9A6", x"7A62091F", x"8FA0C0B8", x"0F75F5A2", x"8B879AB0",
									 -- x"BED98263", x"B1ABC997", x"855580BC", x"BBA8958E", x"7A7B7A78", x"7776787A", x"76716C69", x"6767696D",
									 -- x"6A696765", x"63605C5A", x"5C565355", x"544E4C4E", x"4D4D4A43", x"4141537C", x"93A1A799", x"8C8B816D",
									 -- x"524C7165", x"7BA2CE9E", x"9BAFA27A", x"5D411C36", x"6C90B4B4", x"ABA7998F", x"86A6A4A5", x"96ABA1A3",
									 -- x"85653F2E", x"323C3C37", x"39363430", x"4D92AD8D", x"BA9F5790", x"9B611F14", x"484A565B", x"82715344",
									 -- x"3F578172", x"45643422", x"51440F3A", x"ACC20D5B", x"BA4839B1", x"255E523F", x"97A47479", x"ADB592B1",
									 -- x"7A255083", x"8C8A97A2", x"ABB9B69D", x"9067659B", x"90786869", x"757B8299", x"999490A2", x"7F4AAC8E",
									 -- x"DDDEE2E7", x"E9E8E6E6", x"E7E8EAEB", x"EAE9E9EB", x"EAEDEDEA", x"E9ECEEED", x"EBEDEEEE", x"EDEDEFF1",
									 -- x"F1F0EFF0", x"F2F2F2F1", x"F0F2F5F4", x"F2F1F3F5", x"F2F5F6F5", x"F4F5F4F3", x"F2F4F6F4", x"F3F4F7F8",
									 -- x"F9F8F8F7", x"F7F6F6F6", x"F6F7F8F8", x"F8F8F8F8", x"F8F9FBFD", x"FFFFFFFF", x"FEFFFFFF", x"FFFEFDFD",
									 -- x"FEFCF9F5", x"F1EEECEB", x"EEEEEDEC", x"ECEBEAEA", x"EAEBECEC", x"ECEBEBEB", x"ECEDEEEE", x"EDEDEDEE",
									 -- x"EDECEBEA", x"E8E4DFDC", x"C9C1C1C1", x"B8B4B1AA", x"A9A19F9E", x"9A9DA09C", x"9FA0A3A1", x"9D9EA09D",
									 -- x"A19D9B9C", x"9B999A9D", x"9FA3A6A7", x"A9AEB3B5", x"B9BEC6CA", x"C7C6CBD3", x"D4D7D4D2", x"D9DFDFDE",
									 -- x"DBD6D0C6", x"BFC1BEB5", x"AFAAA39E", x"9C9C9FA3", x"9EA4ABB0", x"B6B9B9B6", x"BAB9B8B9", x"B8B3B1B1",
									 -- x"86677269", x"78716E60", x"6F817A6C", x"4C2330A6", x"5B4E6555", x"407E9D98", x"9C9BAE9F", x"734E5931",
									 -- x"0717150A", x"0F0F3E46", x"4970455A", x"8571463F", x"78465380", x"7D797389", x"7C7C917C", x"7A6F8A86",
									 -- x"69773379", x"8B796775", x"7A735674", x"7A677A69", x"68760012", x"1B296233", x"00131C6D", x"79787C69",
									 -- x"547E8179", x"85838E6A", x"80847F90", x"979B968F", x"7D8C532D", x"88330C28", x"4A468A96", x"76905D6D",
									 -- x"A3216F66", x"A6B2B8AE", x"B19806A7", x"ACAC8EB3", x"AC94B69E", x"92AAB1AF", x"B5CB489F", x"89905704",
									 -- x"036C89A3", x"916F4F9A", x"88687CA4", x"A39E98AC", x"A3B8B1A0", x"838A5335", x"372D60A2", x"AF833810",
									 -- x"2C30466F", x"86A89DA9", x"AD839C9D", x"A5B6ACC1", x"C0B1B360", x"BFDCA3B9", x"A596618A", x"BA9ABDB2",
									 -- x"C2B8DD9D", x"877F5A2F", x"5A8AB097", x"B1D5CFCA", x"CCB39691", x"7E817C80", x"797E7A73", x"747D7371",
									 -- x"6C6D6B69", x"68626564", x"5B625354", x"5659574C", x"47496571", x"879CA3B3", x"C0946994", x"7F835891",
									 -- x"5D769F92", x"A98C7667", x"8B7A5E47", x"0A2F72B5", x"B39DA27B", x"727E879D", x"BB998F98", x"B5B1ABB6",
									 -- x"BEB0C096", x"4B333635", x"39373436", x"6A555846", x"74B39B24", x"8AA06E1D", x"0D3B4D48", x"717A6C75",
									 -- x"A597A3A9", x"4C81A447", x"0D5DB383", x"62657A38", x"52D33C0C", x"953C775B", x"459BA18B", x"9E9C8F9E",
									 -- x"B88E1B05", x"2C7399B6", x"94757798", x"C3B67561", x"5D7E7A8B", x"6E4B6089", x"89918878", x"6C3F7E78",
									 -- x"DDDDE0E5", x"E8E8E8E8", x"E9E8E7E7", x"E7E7E8E9", x"EAECEDEB", x"EBECEEEE", x"EDEEEFEE", x"EDEDEFF0",
									 -- x"F0EFEFF0", x"F1F2F1F1", x"F1F2F4F4", x"F3F3F4F5", x"F2F5F5F4", x"F4F4F4F3", x"F2F4F5F3", x"F3F6F9FA",
									 -- x"F9F8F8F7", x"F6F6F6F5", x"F6F7F8F9", x"F9FAFAFB", x"FAFBFCFD", x"FEFFFFFF", x"FEFFFFFF", x"FFFFFFFF",
									 -- x"FDFBF7F3", x"F0EFEDED", x"EEEEEEED", x"ECEAE9E8", x"ECEAE9E8", x"E9E9E9EA", x"EAEBEBEB", x"EAEAEAEA",
									 -- x"EEEDEBEA", x"E7E4DFDC", x"D6CDCAC7", x"BEB7B0A6", x"A29E9D9C", x"9A9D9F9E", x"A3A09F9C", x"9A9EA09D",
									 -- x"9E999390", x"8E8D8F91", x"91969FA7", x"ABAEB1B4", x"BABBC0C4", x"C1BDC3CD", x"D0D4D4D5", x"DCE0E1E3",
									 -- x"DED9D0C4", x"BAB9B5AB", x"A6A09A97", x"95959799", x"9A9FA4A9", x"ADB1B2B2", x"B3B1B1B1", x"AFAAA8A8",
									 -- x"7C416966", x"606C6E6D", x"98604129", x"010E4A31", x"0B153328", x"3C70877D", x"764F6475", x"818B935E",
									 -- x"4561524A", x"A988677C", x"5B516D31", x"487F7A84", x"4C329277", x"7A765058", x"7D61705C", x"9586726A",
									 -- x"63864951", x"79684571", x"74568574", x"748A6C72", x"5D6B0A01", x"02010004", x"06124575", x"69696869",
									 -- x"5A8A926D", x"98848575", x"71928193", x"918F9885", x"95921458", x"B3AC7332", x"19160505", x"10666AA7",
									 -- x"C55064B7", x"9B8B92D0", x"C45942A4", x"9E97AC9F", x"98BD9FAC", x"B5C4A0CE", x"965880B5", x"DFA8A18B",
									 -- x"5A775F7F", x"98C08553", x"7B480D88", x"9D9A8896", x"90A499A8", x"938E8A95", x"7D4A2955", x"7E807551",
									 -- x"6929255A", x"637C8E93", x"A1A4B9A9", x"8176A397", x"859CDD96", x"50C1C7AE", x"BFC6D435", x"6AB1B1D0",
									 -- x"C1C3ACB6", x"311D58B6", x"DBD1D3B5", x"91ACB2DC", x"DBD9D8CA", x"9F889797", x"A89C9984", x"7574716D",
									 -- x"7076687A", x"6C646464", x"655B6164", x"584C506A", x"8385A6AF", x"9B938C7B", x"827A8A89", x"82968345",
									 -- x"957A5459", x"515F677C", x"52453953", x"968EBCA2", x"6D702B24", x"77908EB7", x"83629D96", x"A1989297",
									 -- x"899E8FB3", x"A37A4F3D", x"31384445", x"56201270", x"56529B9B", x"1E908F5F", x"3007091E", x"43A9A4A9",
									 -- x"9E7074AA", x"A4979096", x"9C643927", x"021F72A2", x"3A3DCF80", x"06701278", x"431F5F77", x"8687938F",
									 -- x"92929A72", x"2E63A193", x"65392948", x"84564F6E", x"62746D56", x"66795D41", x"1E021109", x"6E9F7772",
									 -- x"E1E0E2E4", x"E5E4E4E5", x"E6E5E5E6", x"E8E9E9E8", x"E9E9EBEC", x"ECEBECED", x"EEEFEFEE", x"EDEDEFF0",
									 -- x"EFEFEFEF", x"F0F1F1F0", x"F2F2F3F3", x"F3F4F4F4", x"F2F4F5F3", x"F3F4F5F5", x"F5F5F5F3", x"F4F8FBFB",
									 -- x"FAF9F8F8", x"F7F6F5F5", x"F5F6F7F9", x"FAFCFDFE", x"FDFDFDFD", x"FEFFFFFF", x"FFFFFEFE", x"FEFEFEFE",
									 -- x"FBF8F4F0", x"EEEDEDED", x"EDEDECEC", x"EAE9E8E7", x"E9E8E7E7", x"E9EBEBEB", x"EAEAEAEA", x"E9E8E9E9",
									 -- x"EAE8E7E7", x"E6E4E0DE", x"DED5CFCC", x"C5BCB3A9", x"A8A9A6A2", x"A1A0A0A3", x"A29E9EA0", x"A4ABAFAC",
									 -- x"A39C9390", x"94989692", x"8F91959A", x"9FA4ABB1", x"B1B4B5B3", x"B2B6BBC0", x"C4C7C9CD", x"D3D4D5DA",
									 -- x"DDD6CDC1", x"B7B5B0A6", x"A39D9896", x"95959596", x"999DA1A3", x"A5A9ACAD", x"ACAAA8A7", x"A4A09D9D",
									 -- x"A121222B", x"5F6E5E51", x"472B0600", x"398B5342", x"7497725E", x"02114268", x"667F6876", x"8381926E",
									 -- x"885F6050", x"889B6A82", x"5C70938D", x"6C848A5F", x"5C998C51", x"516B6B62", x"9780767B", x"7C826256",
									 -- x"4F2F3A60", x"9561615C", x"6C687575", x"45505A66", x"7840021C", x"00050200", x"030B334A", x"78757556",
									 -- x"707F7772", x"6C877A67", x"8B7F778D", x"7872917A", x"8B6C0B95", x"9B796683", x"97BEC161", x"050026AE",
									 -- x"85B78C95", x"A3B6BBB2", x"94337BAC", x"5D859E9A", x"9F8EAAAE", x"B0BFBC81", x"58B7B5C6", x"C2BBA5B7",
									 -- x"AE4B0639", x"839892A0", x"D36A008A", x"A7A79FA7", x"A2A5A3B5", x"9FA7A893", x"98A29283", x"6B886358",
									 -- x"804A1B41", x"4456837F", x"9C9EB095", x"92948D80", x"7789A2C0", x"85219288", x"9A89ADCE", x"491C859D",
									 -- x"9F8FB2C1", x"783B89C4", x"C4C3C3B2", x"B4A7ABB2", x"BCB2A1C0", x"BFC8D2E4", x"D9DBD6E0", x"BB9C8B71",
									 -- x"6965746B", x"75657264", x"635F5D60", x"6F8FB58C", x"83AC9A8D", x"7474A3A6", x"B4AFA390", x"86553E41",
									 -- x"512D7196", x"443F6D2B", x"262F5FAD", x"91625A40", x"20627873", x"84848F80", x"70A47C93", x"93676A46",
									 -- x"372E424B", x"73475469", x"6359413D", x"A9B61F1A", x"6154649C", x"89138889", x"566E324F", x"59848479",
									 -- x"86877A9E", x"8D84B26B", x"41423503", x"3E200835", x"2703099C", x"580F390C", x"3A472138", x"6092A282",
									 -- x"7A8871B4", x"8F6AB79C", x"82B0411C", x"040D0500", x"26554544", x"56410002", x"040A0305", x"1C657763",
									 -- x"E2E1E2E3", x"E3E1E1E2", x"E1E5EAEE", x"F0F1EFED", x"E8E7E9ED", x"EEEBEBEE", x"EDEEEDED", x"ECEDEFF0",
									 -- x"EFEFEFEF", x"F0F0F0F0", x"F2F1F0F1", x"F3F4F4F3", x"F2F4F4F3", x"F3F5F7F7", x"F9F9F7F5", x"F6FAFBFB",
									 -- x"FBFAFAF9", x"F8F6F5F5", x"F5F5F6F8", x"FAFCFEFE", x"FEFDFDFC", x"FDFEFFFF", x"FFFEFEFE", x"FEFDFCFB",
									 -- x"F8F5F1EE", x"ECECEBEA", x"ECECEBEA", x"EAE9E8E8", x"E6E8E9E9", x"E9EBEBEB", x"E9EAEAE9", x"E8E7E8E8",
									 -- x"E4E4E4E5", x"E6E5E2E0", x"D9D2CECB", x"C7C1BAB4", x"B8BCB7B0", x"AEAAA8AF", x"B3B0B3B8", x"BDC2C5C2",
									 -- x"B5ACA2A3", x"AFB6AEA0", x"9C9D9B96", x"979DA5A9", x"AAB1B0AA", x"AEBCC1BC", x"C0C1C3C9", x"CFCDCCD0",
									 -- x"D3CDC6BD", x"B6B6B3AB", x"A9A29D9B", x"9C9B9B9B", x"9DA0A3A3", x"A3A5A8A9", x"A9A7A39F", x"9B989696",
									 -- x"958F5213", x"2C2A230C", x"02021D76", x"907A9092", x"7F797874", x"904A1415", x"5B847E7A", x"778A5A23",
									 -- x"6C486F80", x"8B8A976F", x"6B716387", x"9A6F7F93", x"8F747163", x"7262928D", x"70808579", x"607E5B59",
									 -- x"2E588364", x"5851306C", x"653C4567", x"505A656B", x"620E0058", x"7A000202", x"02041324", x"425E9572",
									 -- x"73837E78", x"7B848185", x"868C8862", x"818C965E", x"9B5A0893", x"9B81595A", x"666F7EC3", x"9B603A18",
									 -- x"334A6CA4", x"A1868783", x"6D2E578E", x"64979586", x"949DA5A5", x"A1AF8080", x"C6967FD3", x"ACAEC6A8",
									 -- x"B5A3B774", x"958594BE", x"AFA12656", x"AD909FAF", x"ADB6BAB9", x"AEACA4C2", x"9C8E97A9", x"8B7B9989",
									 -- x"8047622E", x"28353353", x"6E69767C", x"A38DA08B", x"772370A3", x"B0450275", x"A47BACC4", x"AD2D63A1",
									 -- x"8DA3C7D4", x"F16E0FB4", x"BCBA9F73", x"C7A36D93", x"80ADE3B0", x"B4A9767B", x"A2CCC5BE", x"D9DFCEC5",
									 -- x"B691706C", x"717D676E", x"72858D9E", x"9C967B71", x"B1BEB092", x"9BB9A5B3", x"C1919D68", x"4C37322D",
									 -- x"1D46454C", x"6B4D344C", x"7975547B", x"51447091", x"90AC856E", x"9F797768", x"95799CA5", x"8C64312A",
									 -- x"6F99B2B2", x"A7AC888A", x"96BA8D2A", x"11576011", x"0E1F2348", x"B09F5272", x"7F6B6266", x"62338062",
									 -- x"8491A9CB", x"9694A8AB", x"60573C3F", x"4B4B0E18", x"7F620000", x"B9B3543A", x"18322403", x"3264777E",
									 -- x"5C5C7854", x"98969988", x"7590BDB8", x"AC81A48A", x"401C3C15", x"0502101E", x"0E09010D", x"15224967",
									 -- x"DEDEE0E2", x"E2E1E2E4", x"E4ECF4F8", x"F8F9F8F7", x"EBEAECF1", x"F2F0EFF0", x"EEEEEDEC", x"ECECEDEE",
									 -- x"EEEEEEEF", x"EFEFF0F0", x"F1F0EFEF", x"F2F3F3F2", x"F2F4F4F3", x"F4F6F8F9", x"FBFAF9F7", x"F9FCFDFC",
									 -- x"FCFCFBFB", x"F9F8F7F6", x"F5F5F5F7", x"F9FBFCFC", x"FDFCFBFB", x"FBFCFEFF", x"FFFFFFFF", x"FFFDFAF7",
									 -- x"F3F0ECEA", x"E9E9E7E6", x"ECEBEAE8", x"E7E7E6E6", x"E5E8E8E5", x"E4E6E8E9", x"EAEAE9E7", x"E5E4E4E4",
									 -- x"E2E2E3E4", x"E4E2DEDB", x"D1CFCAC7", x"C5C0BDBD", x"BFC3BFB8", x"B7B4B4BD", x"C5C3C5C7", x"C5C6C7C4",
									 -- x"C5BFB8B9", x"C1C6BEB1", x"AAB1B2AB", x"A8AEAFAB", x"AAAAA8A9", x"B2BEC1BD", x"C0C0C1C8", x"CFCDCACD",
									 -- x"CDC8C4BF", x"BABBB9B2", x"AEA8A19F", x"9F9F9E9E", x"9EA1A3A3", x"A3A5A6A5", x"A8A5A09B", x"96949392",
									 -- x"928F9D65", x"1C17040B", x"0C28647D", x"607FA66C", x"7E636F82", x"5F7A8737", x"055A8677", x"778D665D",
									 -- x"8993849D", x"877B5F58", x"66876B92", x"948A8685", x"725F6C69", x"5074807D", x"6A797368", x"6D51575D",
									 -- x"5F888C64", x"3B7B6263", x"4F727F55", x"7A776F5F", x"23000437", x"A7671118", x"0A020008", x"00182F6D",
									 -- x"7F8788A3", x"957C7584", x"8FAA8D9C", x"61929387", x"B0026BA3", x"9D787473", x"85AAAF88", x"A09FC29A",
									 -- x"7C071E22", x"31546E74", x"5C322782", x"97927980", x"838AA48B", x"97B7C0BC", x"745794BB", x"828F7D98",
									 -- x"A27C8FD0", x"053B9B7D", x"789B9705", x"5FAB88AA", x"B4ADBBBD", x"AFA89EA8", x"AAA990A0", x"B7CEAB88",
									 -- x"A7A0704F", x"1E2A2404", x"2D555789", x"9F997878", x"8069467C", x"A4A71054", x"CD95AB87", x"B43A00A5",
									 -- x"D1AA90AC", x"AB825ACC", x"B5DFBDA8", x"BBA7795F", x"525B436D", x"B4AFB6A6", x"6083C0B2", x"BDC6C8C0",
									 -- x"C1D1B287", x"767C8FB3", x"C5C9AA7C", x"79C7B0C3", x"B0A19B88", x"91BA8F91", x"7B326558", x"4C525955",
									 -- x"6B505F87", x"BEB7AFBD", x"C8C9A9B1", x"A2CEB896", x"848F977D", x"88927D7E", x"358AA39F", x"6F202CA1",
									 -- x"BABF9E88", x"9B958F99", x"9286A89E", x"55173037", x"1E00071F", x"92B9C76F", x"58617E5E", x"72674586",
									 -- x"B19DBA81", x"9294A2BE", x"95705867", x"565C9365", x"ABB3A030", x"1EA0E487", x"81372863", x"2E014E99",
									 -- x"9879809A", x"8FB0526E", x"5E56AABE", x"CCB7A1A1", x"958A7163", x"5D4C4B39", x"15180B00", x"0B1A1B3B",
									 -- x"DDDEE0E2", x"E1E0E2E4", x"EAF2F8F8", x"F7F8FAFA", x"F1F0F2F5", x"F6F5F3F3", x"EFEFEEED", x"EDECECEC",
									 -- x"ECEDEDEE", x"EDEDEEEF", x"F0EFEEEF", x"F0F2F2F2", x"F2F4F4F3", x"F4F6F8F8", x"F8FAFAFA", x"FBFDFEFD",
									 -- x"FDFDFCFC", x"FBF9F8F7", x"F6F5F4F5", x"F8FAFBFA", x"FBFAF9F8", x"F8FAFBFC", x"FEFEFFFF", x"FFFEF9F6",
									 -- x"ECE9E4E2", x"E2E2E1E0", x"E6E5E5E3", x"E2E0DFDE", x"DFE1E0DE", x"DFE6EBED", x"EFEEECE8", x"E4E2E1E0",
									 -- x"E0DFDEDD", x"DBD7D2CE", x"CFCEC9C4", x"C3BEBBBF", x"C0C2BFBA", x"B7B5B9BF", x"C4C2C3C2", x"BEBDC1C2",
									 -- x"C7C6C4C3", x"C4C5C5C3", x"BAC3C6C1", x"C0C5C5C0", x"B7ACA9B3", x"BCBCBDC1", x"C1C3C3C9", x"D1D2CFD0",
									 -- x"D2CDCAC7", x"C3C3C1BA", x"B3ADA7A4", x"A2A09F9F", x"9C9FA1A3", x"A4A6A6A4", x"A6A5A19B", x"97959492",
									 -- x"8E88909A", x"6F192232", x"5A817386", x"7B787676", x"75637B76", x"4B6980A5", x"7756686F", x"584A697F",
									 -- x"70767A77", x"7866385D", x"836F9172", x"777A7179", x"6E5D7661", x"6E82924B", x"74574E73", x"5C6A6D46",
									 -- x"5E668167", x"72498F5D", x"5563694A", x"58475463", x"01060C22", x"88514069", x"535D5E62", x"432D1B06",
									 -- x"24566E69", x"7B707C79", x"97527A93", x"4B763F3C", x"201AAAA0", x"8D937590", x"9570B09C", x"8E7F8BBF",
									 -- x"C4AB8E54", x"5A1F0E5D", x"32003076", x"957D687D", x"94977078", x"8F8D7C96", x"828CA787", x"8CB39B94",
									 -- x"AB939088", x"7EA3926C", x"ADC5D183", x"0A7F9FAB", x"B0B9A8A7", x"B5ACACAF", x"A5A3ACA4", x"B3A1989C",
									 -- x"B3B49373", x"82646C41", x"23161505", x"05196F76", x"98995951", x"7BBF3C17", x"B1A0817F", x"B0AE6600",
									 -- x"5CB8BEAA", x"B6A25B8B", x"BFAFBEDD", x"C8D2A778", x"7285A0B2", x"A8DACFD3", x"925F59A6", x"B2B8C8BE",
									 -- x"C7CBC9CE", x"9B97B58C", x"6A7BAEBA", x"C5A8789F", x"6C907C60", x"4E7C8D99", x"7A5A6130", x"85C38C86",
									 -- x"BB96B9C2", x"C6BDBEA2", x"A4A39BA9", x"A285CDBE", x"64606379", x"A381AD69", x"63A16753", x"4365928C",
									 -- x"8E9F9B8F", x"827E6B69", x"65607499", x"996792AB", x"B4763413", x"214B85D7", x"4745ACBA", x"666D779F",
									 -- x"8CA7B0A4", x"8C76808B", x"A5AC4C6B", x"CD83324A", x"57A5BF6D", x"051C61AA", x"AD627033", x"7A2B1E6A",
									 -- x"836A4A6A", x"95A64269", x"5273AEC9", x"ADC1B39A", x"807D5C2F", x"5F525C86", x"785E6656", x"210E3337",
									 -- x"E0E0E1E1", x"E1E0E2E6", x"EFF4F7F4", x"F2F4F6F5", x"F3F4F5F5", x"F5F5F3F0", x"EEEEEEEE", x"EFEEEDED",
									 -- x"EAEBECEC", x"EBEBECED", x"EFEFEEEF", x"F0F1F2F2", x"F3F4F4F3", x"F3F5F6F6", x"F6F9FBFB", x"FBFCFDFC",
									 -- x"FCFCFCFC", x"FBFAF8F7", x"F6F4F3F4", x"F7F9FAF9", x"F9F8F7F6", x"F6F6F8F8", x"F9F9FAFC", x"FEFCF8F5",
									 -- x"EDE8E2DE", x"DDDEDDDC", x"DFE0E1E2", x"E1DEDBDA", x"DADCDCDD", x"E3EDF1F0", x"F1F0EDE9", x"E5E2E0E0",
									 -- x"DDDBD8D5", x"D2CEC9C6", x"CCCCC5C1", x"C3BEBABE", x"C1C0C0BD", x"B6B6BBBD", x"C1BEBEBE", x"BBBBC1C4",
									 -- x"C1C2C3C3", x"C2C2C6CB", x"C5C8CAC9", x"C9CACCCE", x"C8BFBBC1", x"C5C3C3C8", x"C6CACACC", x"D3D5D3D3",
									 -- x"D4D0CECD", x"CAC9C6C0", x"BAB5B0AD", x"A9A5A2A2", x"A1A2A4A6", x"A9ACABA8", x"A6A7A6A2", x"9F9D9A97",
									 -- x"9C8E8F86", x"8F727B58", x"68787579", x"84797F69", x"4C23305F", x"68899481", x"8F94841C", x"15615E39",
									 -- x"596B627E", x"60564459", x"4C737468", x"7B847B7F", x"6C575046", x"869B9047", x"657F9793", x"57886755",
									 -- x"727C6A74", x"67635F4B", x"5C46386E", x"544A5106", x"03110D47", x"672B0945", x"5A537F7F", x"8B885A87",
									 -- x"4A15001D", x"30567684", x"A96C5B7E", x"6D726991", x"4838AB8B", x"8F7E4C77", x"97747D41", x"9EAA94AA",
									 -- x"AAA390B7", x"AA9D5A00", x"001F3811", x"849C816A", x"74796A78", x"6D7E7F7D", x"573B3A8D", x"AB899386",
									 -- x"8A50A38F", x"AFA9CBB7", x"4EAAB9B6", x"654A8383", x"9B9CB1BC", x"A68FA9AC", x"B4A8B4B5", x"AB86252B",
									 -- x"B9B0969E", x"A6868EB8", x"AC4A596D", x"60310D2E", x"44757677", x"5E847A29", x"9E9381AF", x"A8B9A89A",
									 -- x"0024AF94", x"B8D1CA6A", x"7EAFBECC", x"C1B8BDB7", x"8DADAAA3", x"857DBF9B", x"4EAA8EA6", x"A4C0C8C2",
									 -- x"C8B9AFB9", x"D17A5D52", x"4B9A5F68", x"6946816D", x"75929670", x"508B7D7B", x"666D52C5", x"C3BE8A89",
									 -- x"A0A09E9F", x"87938E87", x"72877E98", x"9E8F8C8E", x"A88B6E79", x"55869A72", x"B7AD9886", x"B27D4338",
									 -- x"38415E83", x"8D989799", x"7E83745A", x"73867880", x"7EC1B953", x"0139547F", x"D86117B3", x"AC7A879C",
									 -- x"B6C2B493", x"88797682", x"81A0A379", x"83A76712", x"5D9C9292", x"A4CBA6A1", x"A6BFC970", x"3569231E",
									 -- x"726D6354", x"5D7B8964", x"A1A892CA", x"A5807078", x"7C8893A5", x"8696B7B1", x"A0848572", x"9D381668",
									 -- x"DEDEDFE0", x"E1E2E7EC", x"F2F6F7F4", x"F2F4F4F1", x"F3F5F4F2", x"F2F2EFEA", x"ECEDEEEF", x"F0F1F0EF",
									 -- x"E8E9EAEA", x"E9E9EAEC", x"EFEFEFEF", x"F0F1F2F3", x"F3F5F5F3", x"F2F3F4F3", x"F5F9FDFC", x"FBFAFAFA",
									 -- x"FCFCFCFC", x"FBFAF8F7", x"F6F4F3F4", x"F7F9FAF9", x"F8F7F6F4", x"F4F4F5F5", x"F4F4F5F8", x"FAFAF7F5",
									 -- x"F5EFE6E0", x"DFDFDEDE", x"DCDFE2E5", x"E5E2DFDC", x"DDDEDFE2", x"EBF3F2EC", x"EFEDEBE7", x"E3E0DFDF",
									 -- x"DBD9D5D1", x"CFCCC9C7", x"C7C7C0BE", x"C4C0BBBE", x"C2BFC2C1", x"B9BAC0C0", x"C0BBBABA", x"B5B3B6B7",
									 -- x"C0BDBDC1", x"C3C2C3C5", x"C5C3C6CB", x"C9C3C3C8", x"C8CAC6C0", x"BFC4C5C2", x"C2C8C8C6", x"CACCCACA",
									 -- x"CECACACB", x"C9CAC7C1", x"BFBCB8B4", x"AFA9A5A5", x"A9A9AAAB", x"AFB2B0AC", x"A8AAABA9", x"A7A5A19D",
									 -- x"967F7577", x"696C697A", x"726C6771", x"67543A53", x"71759597", x"7A757671", x"7075707E", x"664B3B5B",
									 -- x"3F535159", x"524D3F51", x"6F6C7378", x"6B716F5F", x"6A66529D", x"687C7D45", x"76C9826B", x"AC5C5275",
									 -- x"42836447", x"75656873", x"6C5E5C46", x"4D590506", x"0C0F226C", x"5A160003", x"0C5B6975", x"5771626C",
									 -- x"7C5B5121", x"28080916", x"6B76A677", x"819A6B57", x"5F4CAF86", x"87728169", x"767A711C", x"94A65FAA",
									 -- x"A9939690", x"87A4AD66", x"51310051", x"725A858F", x"6F657769", x"5D728689", x"84917B6A", x"8D6C7B68",
									 -- x"8072A1BC", x"72BEAFAB", x"CA6C70CF", x"A0546280", x"A694A599", x"9CB5BC9F", x"AAA890AF", x"A79F9D6C",
									 -- x"829B7EBB", x"ACB4B0A6", x"CECDD0D2", x"B6B5651C", x"1E561D5E", x"8B6E9840", x"A9AF9A8E", x"81A191B7",
									 -- x"9F3501AE", x"D0B8DC61", x"6692ADBC", x"ADAABED3", x"B95A5243", x"54687D9C", x"B2CBBFA9", x"B4C5B4B7",
									 -- x"B8B3A7B3", x"B09A6E96", x"6D666889", x"28849C6F", x"81594B49", x"25676842", x"541095CE", x"B4928F72",
									 -- x"7778767F", x"86535475", x"89767588", x"6F50679A", x"9A394C2D", x"002E193F", x"3E56849E", x"C1A4A3A2",
									 -- x"76825771", x"B0A08030", x"66385D9F", x"808D9985", x"417198B5", x"5F1A2249", x"97E15D56", x"C0999D92",
									 -- x"889AA266", x"66857746", x"44829250", x"5B838B9A", x"4D477488", x"9C8EAA8D", x"7D5E7FC3", x"82668127",
									 -- x"2065796F", x"27475C46", x"705F646F", x"7793C1C9", x"C7BDA1A8", x"9F9C879B", x"94BBA794", x"85873A31",
									 -- x"E0DCDADE", x"E1E2E7ED", x"F0F0F0F0", x"F1F3F2EF", x"EFEEEFEE", x"ECEEEEE9", x"ECECEDED", x"EEEEEDEC",
									 -- x"E8E8E8E8", x"E8E8E9E9", x"F0F3EEE8", x"EBEFF1F3", x"F3F5F5F3", x"F0EFF1F3", x"EEF3F7F7", x"F5F7F9FB",
									 -- x"FAF9F9F9", x"F9F9F8F7", x"F4F2F2F3", x"F7F9F9F7", x"F5F4F3F1", x"F1F2F3F3", x"F0F1F2F3", x"F4F6F6F6",
									 -- x"F7F5F1EB", x"E8E6E2DF", x"DEE3EBF0", x"EEE9E6E5", x"E3E4E2EA", x"F4F1EAED", x"E8E7E6E4", x"E2DFDEDE",
									 -- x"DAD6D7D5", x"CBC6C5BE", x"BCB9B8B9", x"B9B8BABD", x"B7B9BCBF", x"BEBBBBBD", x"BBBAB8B5", x"B3B3B5B7",
									 -- x"B8B6B6B8", x"BABBBCBE", x"BFC0C2C2", x"BFBAB9BB", x"BAB9B7B7", x"B7B7B7B6", x"BABDBEBB", x"B9BBBCBC",
									 -- x"BEBEC0C2", x"C3C3C4C4", x"BFBFBDB9", x"B3B1B1B2", x"B5AFB2B4", x"B7B7B0AF", x"B5B0B1B5", x"ADAAA796",
									 -- x"7E796C6F", x"5A454C66", x"6B68625C", x"5452819E", x"7D727E75", x"826B5284", x"73686B5D", x"55541510",
									 -- x"1C49404A", x"58390C4B", x"795E7A70", x"7867746F", x"907C807D", x"86837F6C", x"94755554", x"77628265",
									 -- x"71656451", x"4E5D566C", x"63593C71", x"580E0721", x"001B2862", x"41000211", x"7266566B", x"76998A6D",
									 -- x"7AA19875", x"8D762D35", x"130C0C4B", x"4A4B684C", x"034DAE83", x"8E78748D", x"7B66A386", x"8D9793AC",
									 -- x"96888A8F", x"99989288", x"A5601B41", x"56363276", x"617A827D", x"606B788B", x"806093A6", x"593A4D41",
									 -- x"4D284A76", x"7D9A6687", x"8891568E", x"C6364E81", x"6E716E87", x"8B7B8C86", x"AFB7C8A4", x"A7ACAFC6",
									 -- x"BA9F4A78", x"473C7F75", x"5490ABA0", x"BBC18D54", x"4F818F47", x"8E9F9253", x"79D4A178", x"A9866E27",
									 -- x"D1F8DA24", x"77C09253", x"55698CA6", x"9EB3A8B9", x"A32A3C86", x"A89B9FC9", x"DABAA1B5", x"B7B8C5D1",
									 -- x"C491A0BB", x"AEBA986B", x"76946CB4", x"85756B1B", x"545580A1", x"80A17E7D", x"5A4D3E1D", x"8DA88E5A",
									 -- x"77553C6B", x"9F836E51", x"6A89643F", x"4D615127", x"04203843", x"69534935", x"150E0005", x"1D618492",
									 -- x"BBB1B6A7", x"9097A09F", x"6B666630", x"4EC7B49C", x"94979DB0", x"B3953E01", x"3ABCBC60", x"8A706073",
									 -- x"6A888892", x"B89191A4", x"C76A3840", x"60745E44", x"711B1C29", x"556A6977", x"926A3C9E", x"997D64AD",
									 -- x"674A4277", x"93380101", x"618AACD4", x"CFD56F8B", x"A7AA9AB2", x"A79A949F", x"9D8CB0A5", x"A9A37745",
									 -- x"DDE0E1E1", x"E2E6E9E9", x"E6E9ECEE", x"F0F0EDE9", x"E9E7E7E8", x"E9EFF4F1", x"EAE7E5E6", x"E7E9E8E7",
									 -- x"E7E8E8E8", x"E9E9EAEB", x"EAECE8E5", x"EBF2F3F4", x"F3F3F3F1", x"EFEEEDED", x"F0F3F6F6", x"F6F7F8F8",
									 -- x"FAFAFAF9", x"F8F6F4F2", x"F0F1F2F5", x"F7F8F6F5", x"F1F0EEED", x"EDEEEFEE", x"EFEFF0F1", x"F3F4F4F3",
									 -- x"F0F2F4F3", x"F0EADFD6", x"E1E6EAE8", x"E5E5E4E2", x"E5ECF0F3", x"F7EEE6EA", x"E4E3E2E3", x"E2E0DDDB",
									 -- x"DCD8D5D1", x"C9C4C0BB", x"B9B5B2B2", x"B2B2B3B5", x"B7B5B5B7", x"B9BABEC1", x"B9B8B7B3", x"B0AEAEAF",
									 -- x"B1AFAFB1", x"B2B3B5B7", x"B6B7BABA", x"B6B0AEAE", x"B1AFAEAD", x"AEAFB0B0", x"AEB0B2B3", x"B3B5B6B5",
									 -- x"B7B8BABC", x"BCBBBABA", x"B7B6B6B8", x"BBBBB8B5", x"B9B5B9B9", x"B9B9B4B6", x"B6B5B1AB", x"ADB19D76",
									 -- x"83746F58", x"50625665", x"703F4B6D", x"75826677", x"74714E5B", x"677D8B78", x"5B676B58", x"51461A17",
									 -- x"0000221F", x"3A112B47", x"7C857165", x"875D6082", x"7E8EA78F", x"A38E7981", x"78768977", x"6A90654F",
									 -- x"6C839F73", x"6F776E84", x"625E6A6A", x"281E831A", x"03143E4B", x"59491466", x"44324261", x"68787E62",
									 -- x"82627691", x"94777891", x"75664328", x"15106443", x"309AAC3D", x"5F7E648F", x"B173A87C", x"97AE9A8B",
									 -- x"78553F95", x"738198A6", x"89894D5B", x"30393502", x"3E70746E", x"5A569BC7", x"A193FD8E", x"4B35505B",
									 -- x"5972716D", x"7B6D7E59", x"60897898", x"B516549A", x"014E418D", x"8F919FBF", x"ACA5BCB9", x"B9ACAD89",
									 -- x"AAB9CDC8", x"782E182A", x"331F263A", x"7BB4B5A5", x"81404130", x"506F9253", x"58B39C95", x"A5A1B433",
									 -- x"8BAF9E30", x"14A58493", x"70268788", x"95B5440B", x"45A2C0BB", x"CD9BC7CB", x"C8D2D6C0", x"C1D5D7D5",
									 -- x"E1C68B93", x"A1A89D8C", x"8FA0898F", x"B2923547", x"937C96BC", x"92607742", x"187A4922", x"1F4D6032",
									 -- x"2630232C", x"030E0C09", x"00020000", x"02082253", x"7AB2BCBB", x"C3A8AACE", x"AFA89B72", x"51271C10",
									 -- x"004C5571", x"B1A05252", x"BF3F8BB4", x"BBB1B2CF", x"AEAC9960", x"67B79762", x"28456455", x"6A636777",
									 -- x"888B7DA6", x"AA756E88", x"571A5EA6", x"9D909642", x"80840657", x"3C054D83", x"85836E7A", x"92A2755D",
									 -- x"BEAB80A2", x"8E6D7FA6", x"746CC9B1", x"A2DCA29C", x"ABA89CA1", x"A8ABB8B2", x"A07791AC", x"A399751B",
									 -- x"DAD8DADD", x"DEDDE0E5", x"E6E8E9E8", x"E9EAEAE9", x"E8E4E4E7", x"EBF2F6F2", x"EDE8E4E2", x"E5E7E7E5",
									 -- x"E7E7E8E9", x"EAECEDEE", x"EEEEE9E7", x"EFF5F4F2", x"F5F4F3F3", x"F3F3F1EF", x"F5F6F7F7", x"F8FAF9F8",
									 -- x"FAFAFAFA", x"F9F6F3F0", x"F0F1F3F4", x"F5F5F4F3", x"F1EFEDED", x"EDEEEDED", x"EFEFEFF0", x"F2F2F2F1",
									 -- x"F1F2F3F2", x"F1EDE4DB", x"DEE8E9DB", x"CFD1DDE5", x"EAF3F4F4", x"F5ECE3E4", x"E6E4E2E1", x"E0DFDBD8",
									 -- x"D8D6CFC9", x"C6C0BAB8", x"B7B3B1B1", x"B2B2B1B1", x"B0AEAFB3", x"B6B6B5B4", x"B5B5B4B1", x"ADABA9A8",
									 -- x"AAA9A9AA", x"A9AAACB0", x"ABACAEAF", x"ADA9A9AB", x"ACABA9A9", x"AAACAEAF", x"ABABAEB0", x"B1B0AFB0",
									 -- x"B2B5B7B7", x"B6B4B3B2", x"B3B3B7BD", x"C2C3BFBB", x"B9B7BBB8", x"B6B6B3B8", x"B3B9B0B4", x"B9917182",
									 -- x"71646A63", x"657E778B", x"5573AB9B", x"8B6F6484", x"706D4863", x"5E728A6F", x"49466162", x"5245423A",
									 -- x"6E401C16", x"00107325", x"61785C53", x"3B455A86", x"837B79A8", x"8F7F917E", x"75676985", x"8096468C",
									 -- x"915A766C", x"6D6E6B6E", x"5C745D35", x"0C472908", x"092B6882", x"75667674", x"75783D41", x"94386F44",
									 -- x"64767D74", x"88808CA1", x"94579184", x"7B2A001D", x"5B737F85", x"8AA78E6F", x"75735C7B", x"93817EA5",
									 -- x"6F999478", x"7C8194A3", x"A0913A85", x"93574134", x"1A1E3441", x"4C76A6B2", x"A87D5325", x"58B0CEC3",
									 -- x"BBC3AD7F", x"677D7874", x"7EE1D4CE", x"2283A8A5", x"6E366AAC", x"AD989D71", x"9EC29FAF", x"A59FACAA",
									 -- x"B5C7BAC3", x"C2C3B86F", x"8156372D", x"44338195", x"B69A586A", x"3C5F9878", x"98C39D9A", x"B8E4AA41",
									 -- x"64A55CCD", x"2166F1AF", x"D0301398", x"9A4F0D82", x"CEC3CDB3", x"BEC3BCCD", x"BDC6CACB", x"D7C4C4CD",
									 -- x"BCCBB6A0", x"8D918B82", x"7F8E8687", x"5D5581A7", x"9E565E92", x"84403643", x"90C8D0A8", x"690A3A90",
									 -- x"495C5843", x"60636A5D", x"53705D3A", x"6A8376B6", x"A2939083", x"96A89E97", x"7AB6A6A3", x"D4CBC4A3",
									 -- x"93762D1D", x"004B7C70", x"81B8978E", x"9BA4969B", x"ADB4A66A", x"6990728C", x"A45A013D", x"344C6F83",
									 -- x"934F536B", x"514A323E", x"6F97645E", x"939D8478", x"45858C23", x"3843263F", x"72965F5E", x"81B7D9A0",
									 -- x"7A94B7A6", x"8F8CA2B9", x"9E4841AB", x"B89BB2B5", x"99ABA79D", x"A3AB91B6", x"B4B6959D", x"B9908A89",
									 -- x"CBCDD2DA", x"DFE2E5E8", x"E6E9EAE6", x"E3E2E4E5", x"E8E5E7EE", x"F2F7F6F0", x"EFEBE6E3", x"E4E5E5E5",
									 -- x"E4E5E6E8", x"E9EBEDEE", x"F1F1ECEB", x"F2F6F4F3", x"F4F4F4F5", x"F7F8F8F8", x"F8F9F9F8", x"F9FBFBFA",
									 -- x"FAFAFBFB", x"FBF9F6F4", x"F4F3F1F1", x"F2F2F3F2", x"F1EFEDED", x"EEEEEDED", x"EDECECED", x"ECECEDEE",
									 -- x"F1EFEDEC", x"EDECE8E3", x"DBE2E2D6", x"C9C8D2DC", x"D8DCDADE", x"EBEFEAEB", x"EAE9E7E4", x"E3E2DFDD",
									 -- x"D7D5CAC2", x"C2BCB4B3", x"ADABABAD", x"AFAEABA8", x"A7A8ABAE", x"B0AEABA8", x"ACACAAA9", x"A6A4A3A2",
									 -- x"A0A0A1A1", x"9F9EA0A4", x"A3A2A2A2", x"A1A2A5A9", x"AAA9A7A7", x"A8A9AAAB", x"AAAAACAF", x"AFACADAF",
									 -- x"AFB2B4B3", x"B2B2B2B3", x"B5B9BFC2", x"C2C0BFBD", x"B6B3B6B3", x"B0B0ADB2", x"B5ADB4AF", x"96827671",
									 -- x"6F685760", x"5C5D6160", x"9899756C", x"545A6140", x"80837459", x"75975242", x"5E5D5B70", x"603B6C4F",
									 -- x"4B8B7234", x"34616618", x"5B455C52", x"49336A6D", x"96565398", x"617F946C", x"977B4F5D", x"6D663C86",
									 -- x"824E5A70", x"4E98934F", x"8D717012", x"25390008", x"0E40796B", x"306B6B6E", x"66555A56", x"4525637F",
									 -- x"695F7C89", x"8283928E", x"8B739B83", x"91A25E15", x"2C1F2A1C", x"4D7A4752", x"4A697B86", x"8785827D",
									 -- x"8E807A79", x"95787A93", x"67762B78", x"757E6875", x"3D1E4D81", x"6F644F6D", x"4675DAE3", x"CD9D95B0",
									 -- x"8C767E43", x"4C408C8D", x"67664A50", x"9CE0D4A2", x"CE674561", x"74739593", x"8196ADB1", x"A9C0B9CB",
									 -- x"C3BFB7CB", x"B4B69C79", x"C1B48A7F", x"72503E6A", x"6C8F6472", x"713E4F4E", x"705E9D89", x"7AB876AC",
									 -- x"70ACDCD7", x"9F3F4F68", x"3D932380", x"7786CEC6", x"B5AF94AA", x"B6B2B3C5", x"B6B7C9B2", x"B2AA9CCB",
									 -- x"C4C7CCDA", x"DDA87051", x"97A29A60", x"27729295", x"7B826D6E", x"5B449FB9", x"C59EA043", x"10267EBF",
									 -- x"A9BA9499", x"BCB7CB99", x"4D956A53", x"A1764F7F", x"8B90A58A", x"91AD898B", x"908F788E", x"A9829EC7",
									 -- x"AEE2E4A4", x"A1ACC27F", x"72A3896A", x"6D889482", x"8A9290A3", x"A9A5AC91", x"7FAA9E34", x"40485C5A",
									 -- x"5979788D", x"9EA0AFB6", x"B6AA8497", x"8B88909D", x"986D8676", x"3484894D", x"528199A8", x"9D7B6942",
									 -- x"3DBEBE9E", x"A59AAA9D", x"6D8F4573", x"779B9B98", x"88B4A5A5", x"AEAEA19E", x"9E8F6B65", x"775D868A",
									 -- x"B8BFC5C9", x"D1DBE1E0", x"E4ECF1EF", x"E8E3E2E1", x"E5E2E7EF", x"F5F8F6EF", x"E6E5E3E1", x"DFDFE0E2",
									 -- x"E1E1E2E4", x"E6E8E9EA", x"EAECEAEB", x"F1F4F4F6", x"F3F3F4F4", x"F4F6F8FA", x"F7F9F9F7", x"F7F9FBFC",
									 -- x"FDFDFCFC", x"FBF9F7F5", x"F3F1EFEF", x"F1F2F2F0", x"EEECEBEC", x"EBE9E9EB", x"E7E7E7E7", x"E5E3E6EA",
									 -- x"E7E8E9EA", x"EBEAE5DF", x"DCD7D5D7", x"D7D2CCCA", x"C0C0BCC0", x"CED5D5D9", x"E9ECEDEB", x"E9E7E3DF",
									 -- x"D8D2C2B6", x"B5B1AAAB", x"A6A4A3A4", x"A6A6A4A0", x"A0A1A2A3", x"A4A5A6A6", x"A09E9C9B", x"99989897",
									 -- x"92929494", x"92909193", x"98969595", x"9495999D", x"A3A2A0A0", x"A0A09F9F", x"9FA1A3A5", x"A4A4A7AC",
									 -- x"AAACADAD", x"AFB4B8BA", x"BABCBFC1", x"C0BEBCBB", x"B5B0B1AE", x"ADADAAAD", x"ADADAB8D", x"767C7564",
									 -- x"63796351", x"3843696A", x"636C4C59", x"5F636461", x"707E6262", x"5F72736C", x"736B634F", x"4C2F5259",
									 -- x"1E88745F", x"5D752141", x"63798357", x"5548737F", x"40848282", x"746F6782", x"7F729873", x"5F546A6F",
									 -- x"798B7F72", x"70706C68", x"678B4906", x"1B0F0607", x"171C3657", x"7B7C6B61", x"4A525A8B", x"7B767A91",
									 -- x"7C899583", x"7D958171", x"89958B8F", x"9187766F", x"7D593F53", x"3E013135", x"3DCABD42", x"4D73787A",
									 -- x"77857165", x"644C6650", x"5293366E", x"7F8DC298", x"87421C62", x"BAD79C88", x"C9CCDBCB", x"7F967582",
									 -- x"7F6C85C7", x"BF77C2C6", x"A8977BB4", x"D0AFB78B", x"846B683D", x"635C6359", x"7D75869A", x"9E9CA89D",
									 -- x"A9A8B2BD", x"8F786AAC", x"C7C1BBB6", x"A2C2BEC3", x"ABBE812F", x"5E957C3F", x"836F7B92", x"816F90DD",
									 -- x"63AAD09C", x"D5F17200", x"1B0B8CFE", x"C7B176A1", x"A7ABA2AE", x"B8B0A9B7", x"B5BEB1B4", x"C2C0B6C6",
									 -- x"EAD2C4D0", x"CFA2A766", x"388B6A2B", x"86865B7E", x"8E8B6670", x"7B8D70A1", x"A5A9AB43", x"0A488592",
									 -- x"AE9F8D68", x"7A797991", x"9E807AB3", x"876B526F", x"7377653C", x"3672675B", x"55848D7C", x"9B8F7CA0",
									 -- x"7465407A", x"65668B90", x"8C8B7F6D", x"69639290", x"88828A7E", x"99AEB197", x"7D719A82", x"1A2B6861",
									 -- x"77B6AA9A", x"86707B92", x"81688AA9", x"9A9EBAB1", x"BCB78C6A", x"73137C66", x"5EB7B29E", x"8F7449BF",
									 -- x"A68FAE8C", x"BBA899AE", x"B395A793", x"615E6B7B", x"572B291A", x"34465B3C", x"55788489", x"8467819A",
									 -- x"D1C4BDC0", x"BFBECBDE", x"F1F7FCF9", x"F3F0F0F1", x"EAE4E5EB", x"EEF0EFEA", x"DDDEDFDD", x"DCDBDDDF",
									 -- x"E0E1E2E3", x"E5E6E8E8", x"E5E9E9E9", x"EEF0F1F5", x"F3F3F2F1", x"F0F1F3F5", x"F5F8F8F7", x"F6F8FAFC",
									 -- x"FDFCFBF9", x"F8F5F2F0", x"ECEDEEF0", x"F1F0EEEC", x"EBE9E9E9", x"E7E3E3E6", x"E2E2E3E4", x"E2E0E2E7",
									 -- x"E3E6E8E9", x"E9E7E1DC", x"DBD2CFD4", x"D7D2CDCB", x"C7C9C5C3", x"C7C4C5CF", x"E7ECEFEE", x"EAE4DAD0",
									 -- x"CAC1B1A6", x"A4A3A2A3", x"A2A09C9A", x"9A9C9C9A", x"96989A9B", x"9B9C9C9B", x"99979491", x"8F8E8E8D",
									 -- x"8888898A", x"88868789", x"8B8A8B8E", x"8F909295", x"9E9D9B99", x"99989897", x"96999997", x"96989C9E",
									 -- x"A2A5A7A8", x"AEB8BEC0", x"BDBAB9BB", x"BFBFBBB7", x"B0AAABA9", x"AAABA6A8", x"A7A78E71", x"79745D6B",
									 -- x"6067635C", x"5D7E816D", x"705C7758", x"42575457", x"72674D6C", x"8B795084", x"8D677354", x"422F587E",
									 -- x"43344D5B", x"7064415C", x"645B4953", x"39255E49", x"69A09795", x"6E72726B", x"7B647E81", x"8466A051",
									 -- x"6C83916B", x"63578B74", x"6D8D2505", x"0A00040D", x"0F547D87", x"6F6B6964", x"7A556C75", x"7C727A79",
									 -- x"7E829480", x"61857F77", x"7A758987", x"868F887F", x"80ABB894", x"8B99565C", x"2C4B7662", x"6563546A",
									 -- x"6D95697A", x"555D78BB", x"A4B64369", x"889F8381", x"867C500C", x"24759397", x"887A557D", x"80734848",
									 -- x"90C2BAA4", x"A4545D75", x"6AA6E19F", x"A58F6C7F", x"419FBCA0", x"6FB18D99", x"86A5C78B", x"5563A6B3",
									 -- x"AFC0B9B4", x"A198AFB6", x"B6B7B8BB", x"CEA9ADC9", x"B5B6DB83", x"487AA33A", x"79967165", x"4572BAA3",
									 -- x"565365CC", x"CAC8EF7C", x"377C99B2", x"A06E7B6C", x"77B5A7A5", x"B6BEA0AE", x"A9A5B4BF", x"C4C6B0D1",
									 -- x"D2CBC0BD", x"C6889AA7", x"57405154", x"8A9F6383", x"91633D53", x"A26A277F", x"2B3E7C37", x"033D797F",
									 -- x"848D93A9", x"49194877", x"ADAE818A", x"A55E0635", x"434E5A5F", x"613F3200", x"001D1C36", x"1C220607",
									 -- x"19154D8E", x"9D90AF94", x"92938D99", x"999A857C", x"80709483", x"9A9E7564", x"99968256", x"6B211F55",
									 -- x"5D86797B", x"7BA29878", x"3E93B2A1", x"BABFA5BD", x"C3ABB954", x"56322153", x"9AAB9C65", x"53AE957D",
									 -- x"87697D99", x"A3BBA399", x"9E97BBBE", x"AB8A9369", x"536F4A4B", x"917E7A6D", x"809DC5AF", x"5472A79B",
									 -- x"E6D2C6C3", x"B8B1C4E2", x"FFFFFFFC", x"FAFCFEFF", x"F3EBE7E8", x"E7E7E6E3", x"DEDEDEDD", x"DDDDDEDF",
									 -- x"E1E1E2E2", x"E3E4E5E6", x"E6E8E7E8", x"EBECEDF1", x"F0EFEDEC", x"EDEEEEEF", x"F0F2F3F2", x"F3F5F4F3",
									 -- x"F3F3F3F3", x"F2F0EDEA", x"E8ECEFEF", x"ECE9E7E7", x"E8E7E7E7", x"E2DCDCE1", x"DBD9DBE0", x"E1DFDFE1",
									 -- x"E1E4E6E6", x"E4E1DDD9", x"D4D2D1D1", x"D0CED1D6", x"C4C8C8C8", x"C8C2C7D8", x"EBEEEFED", x"EBE3D4C5",
									 -- x"BAB2AAA5", x"A2A3A5A3", x"9E9E9B98", x"97999998", x"93959798", x"9B9C9A97", x"9996928E", x"8C8A8988",
									 -- x"87868586", x"86858789", x"8787898E", x"91939699", x"9C999694", x"94949595", x"9496938E", x"8F939491",
									 -- x"9B9EA1A4", x"ADB7BCBB", x"B9B6B4B5", x"B8B8B2AD", x"A7A3A5A5", x"A6A7A3A5", x"A185796C", x"6F7C6C5B",
									 -- x"5656717A", x"747C5B47", x"88727464", x"568D615D", x"74675D62", x"87797581", x"72536151", x"2513636D",
									 -- x"691B4539", x"3252211C", x"6A635246", x"255A417D", x"89767A7F", x"5F8A7D9C", x"9B798B82", x"7D75705E",
									 -- x"657E8078", x"61708967", x"68510B18", x"0E06001F", x"5588A08F", x"7E7B6557", x"76565F74", x"6C6B867F",
									 -- x"7177887B", x"617B7F78", x"6F6E7E77", x"8D847A71", x"606A5D69", x"40537B91", x"8B874404", x"2A4E7066",
									 -- x"766E472B", x"213A617E", x"596B4E67", x"676180B8", x"8B939962", x"2B324D5C", x"53716C5E", x"5F575FB2",
									 -- x"9C978075", x"8E807F6A", x"3B57787A", x"866E8EBB", x"AA9C9BB3", x"38659867", x"84653284", x"42727E71",
									 -- x"6651646E", x"96BCD2B6", x"BAB1BCB5", x"BFC7B1AF", x"BEBDAEB9", x"A5BCAC4A", x"656F282F", x"64909B81",
									 -- x"5554946F", x"7EC5C0D1", x"61C7DDC7", x"11768A62", x"84A09ABB", x"A7A7ABB7", x"BDBBB2BC", x"C3C3C5C3",
									 -- x"D1CCCEB3", x"B7AAACA3", x"BA524C3C", x"B8D9D3B4", x"B684403B", x"78704454", x"030C3540", x"63A27B9B",
									 -- x"71959F81", x"73464819", x"624B5019", x"3A3A8721", x"98CBA768", x"88708781", x"7F6B4071", x"678984A3",
									 -- x"B9CB9B7D", x"8B7CA630", x"3D857687", x"9D868973", x"7EAA9374", x"66342325", x"4A7F7282", x"4C2D3930",
									 -- x"352E3D38", x"40513492", x"C7A4A09C", x"7B7C7881", x"5F3F2F45", x"8247344D", x"99706342", x"97A78685",
									 -- x"81763640", x"5B635E54", x"6C787D9E", x"89B5BAA4", x"9CC1C2B5", x"B8C9B197", x"808C98B3", x"BFC0A9AE",
									 -- x"F0F8F6E5", x"DAE3F5FF", x"FCFCFBFB", x"FDFFFDFA", x"F7EEEAE9", x"E6E4E4E1", x"E2E1DFDF", x"DFDFDFDF",
									 -- x"DFDFDFDF", x"E0E0E1E1", x"E3E4E3E4", x"E9EAEBEF", x"EAE7E6E7", x"EAECECEA", x"E8E9EAEC", x"EEEFECE8",
									 -- x"E8EAECEE", x"EFEDEAE8", x"E9EDF0ED", x"E5E1E1E4", x"E5E4E5E4", x"DDD5D6DB", x"D3D0D3DA", x"DFDDDADA",
									 -- x"D7DDE4E5", x"E3DDD6D1", x"CFD1D4D5", x"D6D7D6D4", x"D3D4D3D6", x"D7D1D7EB", x"F0F0EEED", x"EEEADACA",
									 -- x"B9B4B4B5", x"B0AFAEA7", x"A6A8A9A7", x"A7A7A6A3", x"99979495", x"9BA3A6A4", x"9895918E", x"8B898785",
									 -- x"89868485", x"8687898B", x"8E8C8C8F", x"9294989C", x"9895918E", x"8E909293", x"90928F8A", x"8D95958D",
									 -- x"95989CA0", x"A8B2B4B0", x"B1B2B2B1", x"AEA9A4A1", x"A19EA2A3", x"A4A5A1A4", x"856F7673", x"6B6E6768",
									 -- x"625A686C", x"63726D6E", x"6F5B6C80", x"66636568", x"71687D47", x"58538D72", x"634D8948", x"22476A7A",
									 -- x"5700254A", x"475D4C31", x"68594957", x"5A536F80", x"57595560", x"817A5A90", x"5D7C77B0", x"87585368",
									 -- x"5F7B805C", x"66505C4C", x"7B38011B", x"00025B85", x"928C978C", x"4E7F4D53", x"605E3477", x"7D768F74",
									 -- x"6A7B777B", x"95978382", x"564E7972", x"7261667A", x"9C48447B", x"765BB455", x"7C84ACBA", x"3D111872",
									 -- x"96916A6D", x"5B446160", x"39735B4C", x"5394AD98", x"8D988DB0", x"6E2B5A94", x"BACAD0B9", x"AAB9A9CB",
									 -- x"CAB19A85", x"A5B88CA3", x"9F67568A", x"BBA2AA98", x"9E968172", x"C6414F9C", x"9E7F7094", x"B5B3B2AD",
									 -- x"B3AECAB2", x"ACA6B6CE", x"C7ACB3BB", x"AF92BEC1", x"B07D8AAD", x"C9C0A325", x"26265B39", x"6A6F719A",
									 -- x"B4628D8B", x"7D8392B5", x"DEBFCBE6", x"2B71CC78", x"92CEB6A5", x"978CC3B0", x"A9A4B4C1", x"C6BCC1C1",
									 -- x"B5CDC9BD", x"B8B0BCA4", x"BB953851", x"ACA8C5C5", x"C5BE8849", x"5A49588C", x"71808F95", x"A1904075",
									 -- x"964A2256", x"A9877072", x"7D455F6F", x"7C593432", x"60672500", x"0004359C", x"5C63AA82", x"618C7C7E",
									 -- x"2B354F4D", x"148A7641", x"6F571B09", x"2E587A7D", x"70615A45", x"1D1C1D1C", x"18152824", x"21332F38",
									 -- x"3E3D3938", x"48393E86", x"6538423C", x"332F3D2E", x"3D47484D", x"38282B48", x"443E207B", x"9E565157",
									 -- x"96A79B92", x"5E676F80", x"785B6858", x"61535C8E", x"999299A5", x"AAAAA7A4", x"A5927354", x"7FA2A691",
									 -- x"F0F5F5F4", x"F7FEFFFC", x"FCFCFBFC", x"FBF5F0F3", x"EFEDEAE9", x"E7E5E2E0", x"E1DFDFE0", x"E2E0DEDE",
									 -- x"DDE0E0DE", x"DFE2E2DF", x"E2E4E4E3", x"E5EAEBE8", x"E9E5E3E5", x"E7E6E2E0", x"DBE1E8EB", x"EBE9E6E3",
									 -- x"E6E7E8E8", x"E8E8E8E7", x"F5F8F7F0", x"EAEAE9E7", x"E5E8EEEC", x"E3DAD1C8", x"CAC7CCDA", x"DFD7CFCD",
									 -- x"CCD1D5D6", x"D6D5D2CF", x"CCD2D4DA", x"D8D3DCE2", x"E3E2E6F0", x"F7F6F2F0", x"F6F8F8F5", x"F2F0E8E0",
									 -- x"CCC8CACF", x"CFC8C6CA", x"CCCDD6DF", x"DCD1CACC", x"B8B6A79D", x"A8B2B1AF", x"ADA59A98", x"988D8890",
									 -- x"8B8B8C8C", x"8D909395", x"92959892", x"96988E95", x"958F9196", x"928E8E8F", x"8F8D8C8C", x"8E8F8E8E",
									 -- x"969A9C9C", x"A1ABB1B3", x"B2AAA4A2", x"A09C9DA1", x"9E9FA19E", x"9CA5A18E", x"746A6D6B", x"5F633E39",
									 -- x"56625B57", x"61686558", x"7E649566", x"61656E8A", x"716A866C", x"65737960", x"666E5D35", x"4175496E",
									 -- x"4B002750", x"4E463E0C", x"434F606E", x"80998B4C", x"5D6D8D67", x"877484AC", x"62617C87", x"737D6659",
									 -- x"6D997162", x"8A856E69", x"6D23190F", x"01597E74", x"817A905A", x"4F9286A4", x"7E736D90", x"8A6A7F62",
									 -- x"496D786F", x"7A799D6B", x"86787876", x"7A779078", x"934B4478", x"4A949EAF", x"806D8FA3", x"86962C15",
									 -- x"1F4E3750", x"56587445", x"3A687F59", x"70929478", x"8F949D9F", x"A6712546", x"9DCECB95", x"7D89AAB3",
									 -- x"B9B79C67", x"93C581AF", x"AB9076B1", x"BC9C8C85", x"9AA7B188", x"7DA8927B", x"83BBA19F", x"A3787F9F",
									 -- x"949C838F", x"80A8ACA9", x"96959997", x"969EB9A1", x"9BB7AEA0", x"8B8EA693", x"727A6164", x"455EB3D2",
									 -- x"D057393E", x"786BB2C8", x"D9CDADA6", x"275DBB6F", x"A9B59582", x"A2B5ABA5", x"AAA2A6A9", x"B5C2C0BD",
									 -- x"C5D1D1C9", x"A9A9CAB3", x"A3ADAC7D", x"A3A6AAB7", x"BBADBFC3", x"A79D86A8", x"A88F968E", x"949E975B",
									 -- x"60680EA2", x"5767A6BE", x"5F010853", x"A17C947B", x"A897842C", x"6C964C29", x"0000034B", x"5372A6C0",
									 -- x"9B387263", x"6393686E", x"ACAEB394", x"3809141A", x"1F253729", x"2F373A48", x"42393C35", x"2F2E2F3E",
									 -- x"3E3D3138", x"40443E36", x"3D474140", x"4742505D", x"553C5C60", x"495B4739", x"3C34518A", x"AF7F798E",
									 -- x"364F7A7B", x"9B5E6DAC", x"906F92A4", x"B0A77D93", x"978397B6", x"B8ACA886", x"7A603B1E", x"0410798B",
									 -- x"E9E8F3F6", x"FCFFF9FC", x"FCFDFBF4", x"ECE9EDF1", x"F1F0EDEA", x"E6E3E1E1", x"E2E1E0E1", x"E0DDDDDF",
									 -- x"DCE1E4E3", x"E1E1E1E1", x"E4E4E4E5", x"E4E3E3E5", x"E7E5E4E3", x"E2DFDAD5", x"D9D8DADE", x"DEDCDDE0",
									 -- x"E5E5E3E1", x"E0E2E5E8", x"F9FEFFFA", x"F7F8F8F6", x"F5F5F9F8", x"F1E9E0D5", x"CDC8C7CB", x"CCC8C6C7",
									 -- x"C6C7C7C8", x"CACAC6C0", x"C9D2D7DD", x"DDDBE4E8", x"E7EDF4FA", x"FDFEFCF9", x"FAFDFCF9", x"F8F7F1EA",
									 -- x"EBE9E8E7", x"E3E3EEFC", x"FCFBFDFF", x"FDF4EFF1", x"E5E2D5CD", x"D0D0CBCC", x"CBCDC8C0", x"BCB8B0AC",
									 -- x"A49E9CA1", x"A4A3A2A3", x"9D9B9D9A", x"9F9F9294", x"93928F8A", x"8C949285", x"89878586", x"888C8F91",
									 -- x"90949596", x"9CA5ABAC", x"A8A19A97", x"95929498", x"9E989A9E", x"9A948877", x"656E6F6D", x"64575574",
									 -- x"4A6C8279", x"726E5F56", x"627B8D5E", x"5A8C8779", x"73893B7E", x"656B578B", x"716A4437", x"68534A74",
									 -- x"4C041974", x"555A480B", x"14312634", x"3F71534E", x"75737378", x"8B8A92B5", x"7A74A294", x"6D766F8C",
									 -- x"766C7E88", x"74947562", x"39080D00", x"047D7C71", x"7E776F46", x"5F7D725A", x"81746265", x"63898572",
									 -- x"524E416C", x"7583887C", x"836F8B80", x"74766382", x"8A481C57", x"66746C8F", x"8C528AB1", x"69A5DDA8",
									 -- x"57261048", x"5D1B7587", x"59826B52", x"6C85898A", x"9E9D9E9F", x"9FAA8834", x"297ECAC3", x"A1A9B8AF",
									 -- x"A7919699", x"A6CC9F70", x"77753742", x"A4B2A38D", x"8D9E93BA", x"5D66B843", x"6A7A7392", x"ACC08255",
									 -- x"7B818272", x"8CB4A9A0", x"8C878A92", x"8C98AF88", x"97AFC0B7", x"C45A2B5F", x"A6625977", x"AAB2A683",
									 -- x"9D3237B0", x"9994AAAF", x"8E847635", x"101AA67C", x"A79B9FA5", x"99919E8F", x"80B7A7B2", x"B7A9AFB3",
									 -- x"B3B1AE81", x"A6ABCBAC", x"8597A5A5", x"B59FB3C6", x"BCC5B8B0", x"87929B9D", x"73929C9E", x"AB6F5E9F",
									 -- x"80987DAB", x"4A134FAC", x"785F6F8D", x"A7674C4E", x"A381455F", x"7C705D44", x"8578400F", x"2F1E142F",
									 -- x"7AAFB9BC", x"9F757E6A", x"9F812E72", x"B2875530", x"323F3330", x"3F3C3A37", x"4946483F", x"3C333E45",
									 -- x"493E3946", x"4146444E", x"40414D4B", x"47554B4E", x"4F586952", x"4B4D453D", x"3A2D2D25", x"50616ABE",
									 -- x"BF79514D", x"61452447", x"6C7B9FA3", x"8B98C4A8", x"B0908186", x"847B4B42", x"4337353B", x"376EA9AE",
									 -- x"ECF2F6F7", x"F8F4F1F2", x"F0EFF1F1", x"F0F3F4EF", x"EEEDEBE7", x"E2E0E0E1", x"E3E3E3E3", x"E1E0E2E5",
									 -- x"E2E2E1DE", x"D9D7DADF", x"E1DFE0E1", x"DEDADEE5", x"E3E6E6E4", x"E2E1DCD7", x"D4CFCFD2", x"D3D2D5DD",
									 -- x"DFDFDEDC", x"DADCE2E7", x"F5FBFFFE", x"FCFDFCFB", x"FFFCFEFE", x"FAF5ECE0", x"CECBC8C9", x"CBCFD5D9",
									 -- x"D4D0CBCA", x"CCCBC4BC", x"CFDAE0E5", x"E4E4ECED", x"E7F2FCFE", x"FEFFFFFE", x"FCFEFDFB", x"FBFBF8F3",
									 -- x"F1F2F5F5", x"F2F1FBFF", x"FFFFFEFD", x"FAF6F4F5", x"FEFBF6F3", x"F2EAE6EB", x"EDF0F0EB", x"E8EDEFEA",
									 -- x"CEC3B5AD", x"ADAEACA9", x"AAA6A4A3", x"A6A39B9F", x"9794928F", x"8C8F928F", x"88868482", x"8385888A",
									 -- x"878A8B8D", x"939B9F9F", x"9E98918E", x"8C8B8E92", x"94969790", x"8C8B7E67", x"6A767B61", x"774F647E",
									 -- x"51455869", x"75716787", x"6C486B70", x"71817174", x"68564F96", x"74737791", x"69522467", x"6A5D6288",
									 -- x"62171A63", x"426A753D", x"02281E12", x"09000027", x"5468716F", x"95979F96", x"71767D7A", x"846F4A76",
									 -- x"5B73648A", x"58715E64", x"2E030E09", x"258E6674", x"74675E54", x"3E6A5F59", x"705E577C", x"70797E80",
									 -- x"5F4E858B", x"667C7B72", x"797C727B", x"82717D77", x"64610020", x"845E756C", x"60615E71", x"8C9CA97C",
									 -- x"A96D6721", x"082F5B7E", x"376B3962", x"68807492", x"A59D9DA0", x"97B6B0B4", x"73396499", x"CAA7A681",
									 -- x"848FB9C0", x"D1C175A6", x"9E735547", x"426D7784", x"707C3444", x"6AB3719C", x"165A6F70", x"616F7979",
									 -- x"78866E84", x"8299978A", x"82808D73", x"74798C83", x"9586A28E", x"A7AF4266", x"81B6D38C", x"51A15E4E",
									 -- x"9B836EA7", x"9AD0CDA8", x"A7909484", x"BB736E4E", x"939CA89C", x"8F868B6B", x"8490ACA6", x"9DACAEA6",
									 -- x"9E8E92C3", x"E1D3B3B4", x"BFD4C7C1", x"73B2C0AD", x"CCC7BAA2", x"D79E9191", x"7A8AAE99", x"2E394D81",
									 -- x"8DBBA6A3", x"7A42A895", x"915F6D82", x"6E25369D", x"857C706D", x"658B8287", x"95AB8AB1", x"9D919260",
									 -- x"1807539F", x"AC957381", x"9F84777F", x"A37E3D24", x"2D3F3E37", x"485D5559", x"6C524738", x"494D5250",
									 -- x"4146353D", x"46353C42", x"3B404753", x"6C4F5E52", x"577F7E37", x"59583239", x"4C402634", x"392B3042",
									 -- x"53616071", x"9796BA9D", x"5E3A777F", x"74746F6F", x"4A524145", x"3E3B4645", x"483B4A5D", x"96C1B99F",
									 -- x"E2F7EEEC", x"E8E1EFEE", x"EEEEF1EE", x"E7E7EDEF", x"ECEAE7E2", x"DEDCDCDD", x"DFDFE0E1", x"E1E0E2E5",
									 -- x"DFDAD5D3", x"D1CFD1D6", x"D1D0D0CF", x"CDCED7E1", x"E3E8EBE8", x"E7E9E6E1", x"D9D5D3D3", x"D2D1D3D7",
									 -- x"D6D7D9D9", x"D7D7DBE0", x"EDF5FCFE", x"FDFEFDFD", x"FDFAFBFC", x"F9F7F0E6", x"D7D8D8DA", x"E0E7ECEE",
									 -- x"E9E4DEDD", x"DEDCD5CE", x"DDE5E7E9", x"E9E9EDE9", x"E7EEF6FA", x"FBFCFDFC", x"FCFCFCFA", x"FBFCFBF9",
									 -- x"F2F2F6FB", x"FDFAF8F9", x"FFFFFEFE", x"FEFEFDFC", x"F9F9F9FA", x"F9F4F3F7", x"F7F1F2F1", x"EBEDF4F4",
									 -- x"F2ECDBC7", x"BFC1BEB4", x"AEACACAD", x"ADAAAAAF", x"A9A29D99", x"918F9497", x"8F8E8D8B", x"88878787",
									 -- x"83838485", x"8B919392", x"948F8B89", x"88878B8F", x"8F8F8A86", x"8D8D6D43", x"545D525E", x"6D5B464F",
									 -- x"4C064173", x"5D6A7A7B", x"7B79777A", x"7D7C7C6F", x"68638279", x"678A7949", x"6868495E", x"2E54606C",
									 -- x"33410E6E", x"59396C45", x"3639886E", x"4F5E3C49", x"1100285F", x"9068757E", x"867C8D79", x"688E5B99",
									 -- x"757C5B7C", x"806B7A4E", x"200B0C00", x"3B8E7487", x"736A6335", x"61765666", x"88817046", x"11688680",
									 -- x"6A6F5873", x"767D6E61", x"737A6582", x"8E757562", x"53510A03", x"776D6764", x"52717FA0", x"8D7A6872",
									 -- x"B4606E8E", x"4414061A", x"4D996162", x"7488999E", x"979C98B2", x"A0A4B7B2", x"9E2D0629", x"5CA5A9AE",
									 -- x"BEC8C58C", x"C19D58C5", x"AA93B1C8", x"9C463043", x"334F5CB0", x"8E836DCD", x"4C67BF73", x"79917EA0",
									 -- x"AD98A895", x"787799A2", x"7D76555F", x"50565A71", x"876FA3B9", x"B563A2C3", x"A9C9ADCA", x"97453694",
									 -- x"8C9C3A5E", x"8C97AEAC", x"D5B9CDBE", x"6974B994", x"A78F8998", x"73786152", x"8A9C9491", x"8A9C9782",
									 -- x"81ADCDC6", x"B6B9C6BF", x"AE93AED9", x"8278DAB6", x"916AACAD", x"A7B1A99A", x"7D976A35", x"3DA499AF",
									 -- x"6280687C", x"7A413D33", x"4A715C42", x"1F76819C", x"8C929187", x"95AA8B73", x"7581949B", x"AA839D82",
									 -- x"7D340317", x"689487AB", x"8E488B68", x"40293E41", x"5049525D", x"57665F4F", x"50485949", x"4444465B",
									 -- x"6B574A4F", x"5695895D", x"50636441", x"485E615B", x"593B615B", x"9576777C", x"3C4B5548", x"4257564B",
									 -- x"50565230", x"51643E6E", x"6E353645", x"4E463E46", x"4D4F5457", x"50645848", x"5474CEA3", x"68768A82",
									 -- x"E2E6DCDE", x"EBECEDF0", x"E9E6E7EB", x"EBEAEBEC", x"EAE7E2DF", x"DDDCDBDA", x"DAD9D8DA", x"DBDAD9D9",
									 -- x"D2CBC7CA", x"CECFCFD0", x"CBCFD1CE", x"CDD3DDE3", x"E7EDEFEB", x"EAECEBE6", x"E6E5E1DA", x"D8D9D9D7",
									 -- x"D8DADCDC", x"D9D6D8DD", x"E4ECF5F9", x"FAFBFCFD", x"FCFAFCFB", x"F8F7F3EB", x"E8E9E9E9", x"ECF0EFEB",
									 -- x"EDEBE9EA", x"EBEAE7E4", x"E5EAE7E8", x"E9E9EBE5", x"EAE8ECF5", x"FAFAFAFD", x"FDFDFCFB", x"FCFDFEFD",
									 -- x"FDFBF9FC", x"FFFFFEFB", x"FAFBFCFE", x"FFFFFEFC", x"FAF9F9F8", x"F6F6F6F5", x"F7F3F5F5", x"EEEEF3F3",
									 -- x"F0F2EFE4", x"D9D1C9C2", x"C8C3BEBD", x"BAB6B7B8", x"B8B4ABA1", x"A0ABACA1", x"9694928F", x"8C898785",
									 -- x"82828182", x"85898988", x"86848382", x"82828588", x"85888885", x"82807F7F", x"6C5D4E58", x"59594B57",
									 -- x"3C2C2F34", x"5D7A6468", x"7F787D86", x"7D9D7E6B", x"765E5874", x"796B6F70", x"72796E3A", x"68747861",
									 -- x"4D42065B", x"83296B37", x"48167152", x"77646188", x"818F500E", x"2355637C", x"777AA163", x"747A6866",
									 -- x"697D6B73", x"66575747", x"0A030104", x"6E83808A", x"6C671671", x"866F715C", x"594D2717", x"677B7A73",
									 -- x"747C6B84", x"8E6F6464", x"63846771", x"6B6B6B58", x"5775070E", x"4F5E8B62", x"6477A097", x"7E68716B",
									 -- x"405D6B65", x"715F6941", x"19145270", x"609C798D", x"918996A0", x"919FA9C1", x"30309982", x"3A1FB3C3",
									 -- x"8FA9BDC3", x"AB516ABF", x"9B9B9F6B", x"89C7AB8C", x"5E84B489", x"7D887193", x"B1209481", x"72828391",
									 -- x"A3939587", x"6B859483", x"92835958", x"613C7AA6", x"8F808883", x"777B9AA4", x"B4A1ABAD", x"C1B76225",
									 -- x"61921040", x"B47389C8", x"C095AEB0", x"119090B8", x"AD909780", x"785F5472", x"8CAAA09D", x"779F9E8E",
									 -- x"B5B9BFBC", x"C0A4BFBC", x"BF72AAC2", x"B76FCDBC", x"425B71BB", x"9D95A78D", x"7F3155C0", x"608DA968",
									 -- x"4B78431F", x"8DBE6455", x"9EC4BBA6", x"A1B5A098", x"AEB09EA9", x"B4A3AA98", x"A0B28C8E", x"A98F7680",
									 -- x"8C7BAD89", x"2A192A3D", x"424F3C34", x"55515A57", x"59775065", x"754F4553", x"56535663", x"5E5A525A",
									 -- x"4F575858", x"4ECE754C", x"5A46A389", x"5955855B", x"75815087", x"706A816A", x"585B755C", x"334C6D56",
									 -- x"4A4B444B", x"675E4C59", x"4A483D51", x"48445651", x"4656473A", x"375D442E", x"83A74F2F", x"35282A3B",
									 -- x"7A7F999B", x"A5AEADD5", x"F2F0E8E3", x"E2DDDADE", x"DDDBD8D8", x"DADCDCDC", x"DAD7D5D6", x"D5D2CFCD",
									 -- x"D1C8C0C0", x"C7CDD1D3", x"D5DCE1DF", x"E0E5E9E9", x"EAEEF0EE", x"EDEEEDEA", x"E9EBE6DE", x"DEE4E7E4",
									 -- x"EAE9E8E7", x"E3DFE1E6", x"E9EFF5F7", x"F6F6F8FB", x"FCFCFDFC", x"F7F5F3ED", x"EEEDECEB", x"EDEDEAE6",
									 -- x"EBEAEBEB", x"EAE8E7E9", x"E7E8E3E6", x"E9E9EBE5", x"E7E2E5F0", x"F7F6F8FD", x"FDFDFCFC", x"FCFDFDFE",
									 -- x"FDFDFCFB", x"FCFEFFFF", x"FCFCFDFF", x"FFFCFBFB", x"FEF9F8F8", x"F5F6F7F2", x"EEF0EFE9", x"E6EEF5F4",
									 -- x"F5F5F9F9", x"EEDFD9DD", x"E4D8C9C6", x"C5CAD4D2", x"D1C8C1BD", x"BABCBAB3", x"A8A39D96", x"918D8986",
									 -- x"807E7C7C", x"7C7D7D7C", x"7A7A7B7B", x"7A7A7C7E", x"787A797B", x"837E6C5F", x"61668268", x"64515954",
									 -- x"51402200", x"06325E83", x"82736A86", x"835D5563", x"78776A6B", x"716A7A62", x"6F493C47", x"9F77605A",
									 -- x"3C7A1B3F", x"775D3549", x"4A1B6482", x"69658982", x"86969F78", x"23244B77", x"6E8E6D71", x"7E777A6C",
									 -- x"6B66716A", x"5E4E4F21", x"0C00001E", x"9B727371", x"6E263D7D", x"81686A6C", x"472F8C79", x"67617E71",
									 -- x"6485A86F", x"6863585F", x"7386753F", x"616A4858", x"6647001E", x"4C487978", x"6F7D6B45", x"73676961",
									 -- x"1A6D778A", x"7A6D4453", x"BA7A4B2E", x"688A736D", x"70989588", x"9C9BB941", x"2BCBA1A5", x"BC793B98",
									 -- x"C985BDA9", x"A09DB39C", x"A0B59276", x"6C949293", x"67828165", x"6D74AA93", x"B367308A", x"7CAC938D",
									 -- x"92695087", x"94857F7D", x"737C6052", x"714E3A58", x"93716C85", x"B1D4A29A", x"95A79A9F", x"B1BF8D83",
									 -- x"81949531", x"90A76277", x"AEAEBB8C", x"09998180", x"8C61917A", x"7A89A899", x"6497A0A0", x"9399A994",
									 -- x"A6C4B1BC", x"BEB6BCC2", x"B4E0C5BA", x"B81F63D7", x"84D7D6D0", x"CFB4ABBB", x"A23F95AD", x"AA7FA5C8",
									 -- x"C29B979A", x"5F53647F", x"9A908DB3", x"9F7B728F", x"9C9F968F", x"7A81A1A5", x"8B8E8986", x"8FA19CA1",
									 -- x"B2B39F75", x"42224250", x"525E5176", x"638A7A76", x"757A5B56", x"5C585D66", x"42574960", x"4B374142",
									 -- x"41425672", x"6228746B", x"80474360", x"5B4D67A7", x"59856568", x"56515455", x"6952402B", x"4A5E4A53",
									 -- x"1B453F2E", x"4D4E6143", x"35434948", x"3B484555", x"42684F49", x"86674C50", x"45475D5F", x"52574D61",
									 -- x"645D5A57", x"6B73636F", x"8BB0C9D1", x"D7D0C6CA", x"CACACBCD", x"CFD1D2D3", x"D3D1CFCD", x"CBC7C5C4",
									 -- x"CEC9C2BE", x"C1CAD3D7", x"DADEE3E7", x"E9EAE9E8", x"EBECEEEF", x"EFEDEAE8", x"E5E5E2E0", x"E2E8ECEB",
									 -- x"F2EEEDED", x"E9E5E6EA", x"F1F3F4F2", x"EFF0F6FB", x"FAF9FAF9", x"F4F3F1EB", x"ECEBEBEC", x"EDEDEDED",
									 -- x"F2F0EEEB", x"E5E0E0E3", x"E5E6E1E4", x"E5E1E3E1", x"DDDDE2EB", x"F0F1F5FB", x"FBFBFCFC", x"FCFCFCFD",
									 -- x"FBFDFFFE", x"FFFFFEFB", x"FAF6F4F5", x"F4F1F3F9", x"FAF0F1F7", x"F5F3F4F2", x"F6F5ECE1", x"E0E4E9ED",
									 -- x"F1EFECE5", x"DAD3D3D7", x"D3CEC3C2", x"C2CCDEDB", x"D5C8C7CE", x"C9BEBABC", x"C0B9AFA6", x"9E968E88",
									 -- x"7D7B7976", x"75747374", x"73757574", x"73727375", x"6A73736F", x"75756B64", x"4B606F62", x"4F445253",
									 -- x"4F729381", x"2F000B13", x"011F3835", x"8383696B", x"6388755A", x"607B6148", x"67625556", x"55705533",
									 -- x"598B3F27", x"7B695B55", x"4401557C", x"726C6F6F", x"64557698", x"986A440E", x"32435983", x"715C524E",
									 -- x"6F86626C", x"64532D04", x"08060416", x"8B707061", x"54047C59", x"3E5F5943", x"4885676F", x"63767881",
									 -- x"9A62506F", x"596F6C69", x"63506267", x"706B7059", x"4F2B0612", x"47596465", x"59666C9E", x"78766A88",
									 -- x"9377AC6B", x"7D751900", x"5A8E6F37", x"22495A4F", x"404C78B2", x"A8850B2F", x"C2A3ACA7", x"B2E39938",
									 -- x"61BDAE9D", x"95BCB59A", x"9F7592BA", x"A89A9B9B", x"908E9493", x"99A1A99B", x"8F660636", x"6E7B7073",
									 -- x"AFA6909B", x"6D855E6A", x"5659634D", x"7A7885B4", x"AAC6DABE", x"A1A8918F", x"8E9B7F9A", x"A9A9C1C2",
									 -- x"CEB7ABD6", x"82C79594", x"8970A65C", x"71ABAA4F", x"545475A6", x"6A8A99B5", x"926FA5AE", x"A299977E",
									 -- x"68A4AB9F", x"ACBEBEA3", x"B0C0BAB1", x"A95B8BAD", x"9E6D467B", x"80C0CBB7", x"91858587", x"A99E8C62",
									 -- x"855366B3", x"8B9D91A5", x"A59A9A95", x"9D9AAA9F", x"ADA88C93", x"958E8968", x"7D9C6F7F", x"848C956C",
									 -- x"4D4C4335", x"3E538056", x"74A06D46", x"3865365A", x"4051695A", x"7C8C5C62", x"6E69413E", x"32354B4F",
									 -- x"464A5C68", x"73585E6D", x"51223055", x"92A55784", x"7D78476C", x"411F2744", x"4B857163", x"69615A59",
									 -- x"7571505A", x"3E597350", x"5E5A4A56", x"59605C4B", x"2C417949", x"43516D56", x"3C4F6D5A", x"5D6E6C74",
									 -- x"79907466", x"6B6A7670", x"4E676E7B", x"A6C1BEBC", x"C0C1C3C2", x"C1C0C0C1", x"C5C4C3C1", x"BEBABABC",
									 -- x"BEC3C6C5", x"C5CBD2D4", x"DDDDE1E9", x"ECEAE9EA", x"ECEBECEE", x"ECE7E2E0", x"E3E1E0E2", x"E4E5E6E7",
									 -- x"E8E6E5E7", x"E6E1E0E3", x"E5E5E4E2", x"E0E3EDF5", x"F7F6F6F6", x"F2F2F0EA", x"EFEEEEF0", x"EFECEEF1",
									 -- x"F9F6F1EC", x"E4DEDEE1", x"E3E3DFE1", x"DDD5D7D7", x"D3DAE3E8", x"EAEDF3F9", x"FCFCFDFE", x"FEFDFEFF",
									 -- x"FEFEFCFB", x"FEFFFBF4", x"F3EBE8E9", x"E8E7EEF9", x"F5E8ECF7", x"F5F0F2F3", x"F1ECE3E1", x"E2D9D8E4",
									 -- x"E8ECE3CE", x"C5CACCC5", x"BDC4C4C0", x"B2AFB8AE", x"AAA5ABBB", x"C9D0CDC5", x"C1BAB1A9", x"A1968A81",
									 -- x"7D7B7976", x"73717172", x"7071716F", x"6C6C6C6D", x"6D6D6A6E", x"72686067", x"6D625E65", x"6A3F5660",
									 -- x"4D8F7C73", x"91887D7B", x"4456713E", x"1C355A41", x"535F6666", x"5A475A7F", x"82546480", x"65775F5D",
									 -- x"613C5523", x"8F517A76", x"3A174563", x"5E6D615D", x"79726569", x"8D7F8F82", x"60521A22", x"23170201",
									 -- x"1F210A15", x"1D2D2D10", x"03000C28", x"8D726360", x"33349664", x"4C7A3B5A", x"83A3456B", x"82636A77",
									 -- x"787A736E", x"7199654D", x"3F77816F", x"6687505E", x"6F6C001B", x"406D7772", x"6B727F9F", x"78754C67",
									 -- x"5C677659", x"A87C687D", x"5431001F", x"13012934", x"82968995", x"7F3351AF", x"9F9F9CA3", x"BBC1D1D4",
									 -- x"94536497", x"BF94B497", x"8A94667C", x"93B1A09B", x"7D9FC49A", x"8693967E", x"745E1218", x"5B736770",
									 -- x"8B8F9A87", x"604F5842", x"50425AAB", x"917A9F9F", x"B2A59696", x"A2A7A994", x"7B8C94AD", x"9B9EB3B2",
									 -- x"A6C1ABA9", x"7089C3A9", x"8F5E471F", x"38208145", x"2B2445A7", x"829EA9B7", x"D6966896", x"8F757885",
									 -- x"868A9299", x"A3B8BEAE", x"B2B6ACA8", x"8F8ED6AC", x"BB9E8C98", x"3F828B96", x"8C5D667F", x"2A938B90",
									 -- x"AAA4C2AF", x"B19FA193", x"A5B9A195", x"A0B3A5A7", x"A3A28875", x"93917766", x"63AA8F83", x"5F5C4546",
									 -- x"6E594F59", x"733E3E56", x"3F482341", x"53628367", x"6386A184", x"95866497", x"9A7D6C67", x"7D8E7057",
									 -- x"5153765B", x"57562A44", x"6161646C", x"58945159", x"6167897E", x"80B85D79", x"6DA7A68B", x"8E8E5E7B",
									 -- x"5C544F73", x"5037525A", x"8B392D67", x"645F7458", x"545C5F61", x"42394B5A", x"524C4558", x"403D4449",
									 -- x"8C828079", x"797A676A", x"70686A5F", x"50BAB8AD", x"B1B0B5B4", x"B4B3B6B3", x"B9B6B5B6", x"B6B4B4B5",
									 -- x"B6BDC3C3", x"C0C4CCD3", x"D5DADEE2", x"E8EDECE7", x"EAE9E8E8", x"E5E0DDDD", x"DDDDDCDE", x"E3E6E3DE",
									 -- x"DFE4E6E0", x"DBD9D7D5", x"D7D8D6D4", x"D8DCE1E7", x"EDE9E9EC", x"EDEAE9EB", x"EAEBEDEE", x"EFEFF0F0",
									 -- x"F2F3F4F4", x"F0EAE4E0", x"E0DEDEDD", x"D9D5D4D6", x"CCDAE7EA", x"E7E7EBF0", x"F8FCFCFB", x"FFFFFCFB",
									 -- x"FCFBFAFB", x"FDFBF6F1", x"E8E8E6E2", x"E0E4F0FA", x"E9E9F3F9", x"F4F1F1ED", x"EFE2DAE3", x"DBD8D5DB",
									 -- x"E8EAECE1", x"D8D8CDBF", x"C1C5C1B3", x"A9A6A4A0", x"9E9DA1A4", x"D9D6D2CB", x"C7C0B2A5", x"9B8E8584",
									 -- x"807C7C7C", x"75717171", x"6F6E6E6E", x"6C696869", x"696E6966", x"7D77525A", x"70816A6D", x"67667D46",
									 -- x"65807476", x"706F7B7B", x"9B959998", x"7141100E", x"2B6D5F60", x"5B676471", x"8B588878", x"646F5C66",
									 -- x"62794831", x"894F657B", x"55560D4E", x"565E6C69", x"6A746D65", x"726E7979", x"8A971372", x"29051668",
									 -- x"717F7351", x"2D0F0100", x"02030242", x"83605E42", x"014E7067", x"5C543876", x"544F7A8D", x"A2966C6B",
									 -- x"73797273", x"73665D68", x"7552313F", x"30383F6E", x"70884515", x"4E748F88", x"77316C6C", x"61709777",
									 -- x"7489486A", x"86738B98", x"97D78E48", x"5C304A53", x"13508466", x"056DB297", x"97838685", x"A0CFBABB",
									 -- x"BCB66B1B", x"539FAA94", x"8B878486", x"879FA2AE", x"95A29794", x"9291878F", x"9E81704C", x"6C80946B",
									 -- x"A3686B8E", x"8A6D4F66", x"6E8A8989", x"7A8C8C92", x"999D9A92", x"909BC6B8", x"9C95B2B2", x"AFA9ACBF",
									 -- x"B4A89D84", x"C38F23B6", x"7A09455D", x"77642331", x"30501830", x"546AA9AC", x"B8D1A06F", x"958C8ABA",
									 -- x"9A758C9A", x"BDB3B2B2", x"A6A08595", x"8B5881AD", x"AFCFDCBA", x"A793457A", x"7F6DB9B9", x"92708E8B",
									 -- x"8C889891", x"A8A8AAA0", x"93B79391", x"8C959D89", x"8B744040", x"43475355", x"4F555446", x"4C44454E",
									 -- x"533B5F5B", x"6066635B", x"5A818E8C", x"9D8E9059", x"565CA289", x"7685729C", x"61445C5C", x"515C6261",
									 -- x"5A576B6B", x"4F63946F", x"667C7E61", x"5A48205A", x"51556D6A", x"5F686BA1", x"7970533B", x"534A4C4C",
									 -- x"2A2B4846", x"4E465050", x"4C4A4D59", x"525D6B6E", x"74695040", x"514B6675", x"796B5C58", x"5D655246",
									 -- x"86998C80", x"8E7B7678", x"70897642", x"626F8DB9", x"AEADB3AE", x"A7ADB4AA", x"B1B1B1B2", x"B1B0B2B5",
									 -- x"B2B7BABA", x"BABEC4C8", x"C9C9CBD1", x"DDE6E3DB", x"D9DADBDB", x"D9D6D6D8", x"D7D9DBDB", x"DBDAD6D0",
									 -- x"D3D6D6D3", x"CFCCCBCA", x"C7CACACA", x"CED0D3D8", x"DDDADADE", x"DEDCDDE1", x"E5E5E6E7", x"E8EAEDEE",
									 -- x"F1F2F4F4", x"F3F0ECEA", x"E6E7E9EC", x"ECEAE9EA", x"E4EBEFED", x"E9E7E9EA", x"F2F6F8FB", x"FFFFFFFF",
									 -- x"FFFFFCFB", x"FBF8F4F0", x"F1F1EFEA", x"E6E8F1FA", x"F1EFF2F4", x"F1EEEEED", x"E7E5E1DD", x"D3D5D5D4",
									 -- x"E0E7E9E9", x"DACAC7BE", x"B4B4B1AB", x"A5A09D9A", x"9698A1A9", x"D4D5D4D0", x"CDC6B9AE", x"A69A9292",
									 -- x"8B878582", x"79737270", x"6D6B6B6B", x"69676667", x"665E765F", x"1E366761", x"6D776E65", x"4F695C67",
									 -- x"93836661", x"7269556E", x"7474986E", x"67618077", x"4D1E5A5A", x"5A79676C", x"73746373", x"766D735F",
									 -- x"5A592A46", x"9862566F", x"5D03344D", x"595A5762", x"69695669", x"6166687E", x"77006BA8", x"8873946B",
									 -- x"60646D85", x"876F5B32", x"12020075", x"85597619", x"2D705F55", x"3D5B636C", x"5F607172", x"7E719173",
									 -- x"6659636F", x"80704225", x"4F4A5448", x"585C7C71", x"6C62661C", x"3B6A6F5F", x"25587D4D", x"725573BA",
									 -- x"64226183", x"994E3044", x"6D857542", x"7D7E6D81", x"7C30315F", x"44A5A5A9", x"A2848B92", x"93ACB1C7",
									 -- x"A489B0A1", x"24399299", x"8696AD9E", x"AD9BAEA7", x"B1A76F5C", x"97868676", x"5B0C1E33", x"5B7F7978",
									 -- x"876D4D59", x"897B729D", x"8A8B9286", x"B5BF7E74", x"93959089", x"7E6B93C6", x"A9ADADA3", x"B0B0AAA8",
									 -- x"B6A5AD91", x"5FB87C42", x"1975AF6C", x"89C1D777", x"69706A27", x"18174CA3", x"C9C9BF9A", x"A7AD6D85",
									 -- x"63836E8B", x"98919794", x"A5999BA5", x"556FBABB", x"AA71B0B9", x"A0C4B072", x"ABAFACC5", x"D8BEADBF",
									 -- x"90648967", x"5F68776C", x"63716554", x"3D4D404B", x"4E59596F", x"544E5554", x"5A4A4445", x"4948433D",
									 -- x"3F4D5C5E", x"6A9C8CAC", x"EFA48461", x"87735655", x"5B4D5D66", x"75604E50", x"68AE5C7F", x"7F465560",
									 -- x"62368EB3", x"797D9F4A", x"261B4049", x"3013371A", x"4BBE7151", x"4D564644", x"5E5C4F42", x"4B50503B",
									 -- x"3E4E4C5C", x"655D5526", x"3439344F", x"48514536", x"5D666459", x"746E7FA5", x"A580806F", x"6F647576",
									 -- x"7899836D", x"50477A64", x"6F7F8565", x"475A585F", x"A0AAABA7", x"A5AAACAF", x"A8A9ABAB", x"A9A9ACB1",
									 -- x"B0B1B2B2", x"B3B7BABB", x"BDBCBBC0", x"CAD2CEC7", x"C6C7CACB", x"C9C7C9CE", x"CED3D7D7", x"D4CEC9C5",
									 -- x"C7C6C5C5", x"C3C0BEBF", x"BCBFBFBF", x"C3C4C4C8", x"CDCBCCCE", x"CFCFD2D6", x"DCDCDDDD", x"DFE3E7EA",
									 -- x"E8E9EBEB", x"EBEAE8E7", x"E7E8ECF1", x"F3F1EFED", x"EEEFEEEC", x"EBEBEBEA", x"EDF0F0F1", x"F2F2F6FF",
									 -- x"FCFCFCFD", x"FCF8F3EF", x"F4F6F5F1", x"ECEDF3F9", x"F4F5F5F6", x"F6F0EAEA", x"E7DED6CB", x"C9CED8D7",
									 -- x"D9E3E3EA", x"D1AEAFAA", x"A7A19E9F", x"9E999593", x"90939BA4", x"BEC4C8C8", x"C4C2BAB3", x"AEA59E9E",
									 -- x"948D8883", x"7973726F", x"6B696766", x"64626162", x"6A635764", x"58371E28", x"384B4B3A", x"5E53255F",
									 -- x"8E756669", x"6E6E5567", x"587E796B", x"4D441489", x"8E431C27", x"4968705A", x"6B78567D", x"8A6F613C",
									 -- x"56553C37", x"7C3F3939", x"5D743920", x"4D5C4537", x"48555A67", x"5E6B6147", x"3E2B7870", x"747C747F",
									 -- x"6E648277", x"7D897E87", x"82725A6C", x"67742F1A", x"86676972", x"6B65736B", x"8A86756B", x"65586147",
									 -- x"716F536A", x"3C00163D", x"70747D67", x"6464844A", x"557F6916", x"17475440", x"2D7E548F", x"6E55481F",
									 -- x"14498D82", x"4B3EA1D6", x"79013831", x"6487512D", x"98C67501", x"3A80A38F", x"8E90859A", x"9CB0CDB5",
									 -- x"BAB29893", x"B086113D", x"66788071", x"93BA8559", x"5A788C89", x"95683D0B", x"00558CB9", x"C4986A79",
									 -- x"A5BC7494", x"674E8180", x"96777D97", x"7B75828E", x"795D79AB", x"AFAAB8AA", x"A4A0AEA1", x"A9B8AA9A",
									 -- x"A9A4A8AE", x"B8B299B1", x"534F4F45", x"37052D68", x"ABCAB15B", x"343E2D2C", x"56A4B8B7", x"81B3AE97",
									 -- x"9D6984A3", x"738DB99A", x"795F8E6E", x"2061CBB0", x"B178818E", x"757D7674", x"B6927F72", x"94ADB2A8",
									 -- x"B0A43D36", x"25262E35", x"444A5A5A", x"55715967", x"76575652", x"47384C4C", x"38435049", x"4A4A5968",
									 -- x"5E665E4F", x"9175A0C6", x"AF696853", x"8A804B5C", x"89634E77", x"78997559", x"5F998499", x"C2896890",
									 -- x"89AA7D5C", x"5D4A4A52", x"81855558", x"554B6567", x"565B2C58", x"56475459", x"59414351", x"4B424431",
									 -- x"4E636456", x"3B386353", x"3F474B64", x"51635162", x"8B727063", x"6C696F82", x"73506869", x"6755645A",
									 -- x"7A65746B", x"648B9782", x"8B81877D", x"767B7554", x"4A91B0A3", x"A6A6A0A6", x"A3A4A5A5", x"A4A4A8AD",
									 -- x"B0B1B0AE", x"AEB0B2B2", x"B2B5B7B8", x"B9BCBDBC", x"BABABCBD", x"BCBBBDC0", x"C2C7CDCE", x"CBC6C2C0",
									 -- x"C0BBB9BB", x"BBB8B6B8", x"B9BBB8B6", x"B9BABBBF", x"C0C0C0C2", x"C2C2C6CC", x"CDCDCECF", x"D1D5DADD",
									 -- x"DCDDDFE1", x"E2E2E2E1", x"E4E6EAEF", x"F2F1EEEB", x"E9E8E7E8", x"EBEDEFEE", x"ECEBE8E5", x"E3E2ECFC",
									 -- x"FDFDFEFE", x"FEFBF8F6", x"F6F8F8F6", x"F6F8FBFC", x"FAFAF4F1", x"F2EBE2E3", x"DABEB1B0", x"BCBDC9CE",
									 -- x"CFD6DBE3", x"CCAAA9A9", x"9E999595", x"95928F8D", x"8D8C9097", x"A2ADB7BA", x"B9BBBAB8", x"B8B2ACAC",
									 -- x"9F958B83", x"7B77746E", x"6C696665", x"64626263", x"5A676768", x"66777472", x"6A746A7C", x"787A8375",
									 -- x"818C6363", x"796C7460", x"685F5563", x"8F835954", x"636F885C", x"05187B95", x"815C5F67", x"63625770",
									 -- x"5850210F", x"2A124063", x"6C665400", x"30373B3C", x"3450614A", x"645D5435", x"146E7B54", x"8C788682",
									 -- x"75797572", x"86746973", x"6A858769", x"47002182", x"9B816A61", x"69706585", x"8C605169", x"605C6A5F",
									 -- x"65402A08", x"044C4E54", x"8777495F", x"646B617B", x"736C4A73", x"3B07581E", x"435A6A7B", x"39584D60",
									 -- x"93B35D6E", x"56797493", x"76594478", x"9284803F", x"525ED57F", x"40234CA7", x"86AC956D", x"7C9EAAAF",
									 -- x"AABA8A66", x"A0B47025", x"000C0A0B", x"111C0A2B", x"37B1AEAF", x"9A8786B0", x"BBC7B1A4", x"92A3A290",
									 -- x"67868690", x"B098688D", x"98795358", x"6C6A8052", x"67576E81", x"7D8A9398", x"97BAA2A8", x"B6A2ABA7",
									 -- x"A8A3AFC1", x"A3B4B8A7", x"B89082B3", x"C887AC7E", x"3F505F75", x"6D86DDAE", x"371E7199", x"825598AE",
									 -- x"9C5C8691", x"9696B580", x"73738B94", x"984B7E9F", x"A0B1D0C0", x"B3B8DABE", x"92B1A99A", x"535F8E88",
									 -- x"7A715151", x"6F7A6C86", x"77756C66", x"656D605A", x"684C4E40", x"64BB593E", x"4C5E665A", x"5E538F8A",
									 -- x"7F976165", x"57465D54", x"525B5F35", x"4F676567", x"7E6E9785", x"7B8A898C", x"7B5E5D4D", x"66C6A762",
									 -- x"525A564D", x"4669494C", x"61646D61", x"4D425660", x"634B3D48", x"595F565E", x"6A5D5C8E", x"5A4D393E",
									 -- x"553E5064", x"87695A64", x"6171755E", x"54916F6A", x"7E5B5D63", x"6C696860", x"635A5D80", x"63745643",
									 -- x"83787C7C", x"9A6E6569", x"87537961", x"7C8D7590", x"685A5559", x"999EA5A5", x"A2A1A1A1", x"A2A3A6AA",
									 -- x"B1B3B2AD", x"A9A8A9A9", x"A7ACAFAF", x"AEB0B3B5", x"B3B1B2B4", x"B5B4B4B5", x"B7BABDC0", x"C0BEBDBC",
									 -- x"BAB4B0B2", x"B3B2B0B1", x"B3B4B1B0", x"B2B3B2B5", x"B6B6B7B7", x"B6B7BBBF", x"BEBEBFC0", x"C1C4C7C9",
									 -- x"C9CACED1", x"D3D5D5D5", x"D7D9DEE3", x"E8EBEAE8", x"E7E5E3E2", x"E4E6EAED", x"EAE9E6E3", x"E1E0EAFB",
									 -- x"FFFFFDFB", x"FBFBFBFB", x"F5F6F5F5", x"F8FBFBF9", x"FEF9EBE2", x"E2DDD9DC", x"C8A89EA5", x"B3AEB5B9",
									 -- x"C2C3CCCC", x"BCA9A1A2", x"9997918B", x"89898886", x"8785868D", x"919FABAF", x"AEB3B4B4", x"B7B5B2B2",
									 -- x"AEA39993", x"8C888278", x"6E6A6563", x"61606061", x"65676364", x"686B5F6C", x"7B687352", x"6D54447B",
									 -- x"61536867", x"6E707778", x"3E38615B", x"6C59608D", x"8C708470", x"60130B47", x"416D6B54", x"48516E53",
									 -- x"5C4A1106", x"383D5C42", x"5B6E5510", x"0D352C30", x"3A4B4635", x"64432528", x"2E575353", x"546A9D7F",
									 -- x"7D85736E", x"725D7AA4", x"9D7B6A62", x"642D2C6E", x"7E706C66", x"5B5F6264", x"5E695862", x"815E4710",
									 -- x"0014597A", x"95A23D5E", x"776B836D", x"5F4E536D", x"5F625A50", x"872D2020", x"6341681E", x"437D2A2B",
									 -- x"819B5026", x"7B662E24", x"AE8F604E", x"AE511A7F", x"856341A4", x"92B59C4B", x"80B09189", x"8594CAA1",
									 -- x"86A69B94", x"9C8AA292", x"927D8B83", x"6D7039A7", x"A589707A", x"6BA3908E", x"91988A93", x"9FA2ADBE",
									 -- x"A282928F", x"8087897F", x"7E957B63", x"5378676C", x"8695738E", x"725F9388", x"889899A7", x"A6A3B6B4",
									 -- x"A89D8582", x"62ADB99F", x"AEABAA7F", x"74D7B7C0", x"B2B0E3B4", x"82B2C3C4", x"E27B245D", x"566B8686",
									 -- x"8A81A393", x"B5807BA0", x"B8C3B0B4", x"7D51B285", x"8994718E", x"94989582", x"5E797173", x"66654D68",
									 -- x"6F584E97", x"C27D6176", x"4F5D6464", x"6554606A", x"5C4D6066", x"69F5A252", x"82786A5B", x"656D3362",
									 -- x"7DB18F76", x"745D6382", x"3C60663E", x"556C7433", x"4A495B42", x"59393330", x"585A4F6C", x"575D995D",
									 -- x"5F545960", x"37464D6B", x"57516C52", x"514D4D61", x"6B657D7D", x"5E807F4B", x"6B666174", x"5C5D5E64",
									 -- x"6E5A6B6A", x"677E818E", x"7385866E", x"6D977961", x"716B5E5F", x"665B6168", x"69585E53", x"5F5A5745",
									 -- x"7981616A", x"655B3D76", x"6864735B", x"46665D7B", x"5C654650", x"52979A97", x"9D9B9B9C", x"9D9FA3A7",
									 -- x"B0B2B1AB", x"A4A09F9F", x"A0A0A1A2", x"A4A5A5A5", x"A9A8A9AD", x"B0B0AFAE", x"B0B0B1B4", x"B5B5B5B5",
									 -- x"B3AEA9A9", x"AAAAAAAA", x"A7AAA9A9", x"ADACAAAB", x"AFAFB0B0", x"B0B1B4B6", x"B7B8B9BA", x"BABBBCBD",
									 -- x"BCBDBFC0", x"C1C1C1C0", x"C5C8CCD0", x"D5D9DBDA", x"DEDBD7D4", x"D3D6DCE1", x"E1E4E3E1", x"E0DEE2EE",
									 -- x"F8F9FCFF", x"FFFFFBF7", x"F7F6F4F3", x"F5F9F7F2", x"ECE6DDD8", x"D7D4D2D4", x"C0ADA3A1", x"A3A2A8A9",
									 -- x"AEACB4AE", x"A29B918E", x"92908B82", x"7E7F7F7C", x"7F7D8086", x"89939C9F", x"A6AAAAA9", x"ACADACAF",
									 -- x"B0AAA7A5", x"A2A09A90", x"847D756F", x"6B676565", x"67697171", x"727E785A", x"74817163", x"41516875",
									 -- x"6F7D4B6B", x"6E84743B", x"78853833", x"30543D4F", x"6A576B62", x"5E726E3B", x"12312F40", x"5748543D",
									 -- x"270B0011", x"39173B3A", x"4D41411B", x"00262631", x"37423832", x"2F443E46", x"1A52554F", x"554B5E53",
									 -- x"474D5859", x"5966696A", x"70566E76", x"25554C08", x"314F886B", x"5D5C5757", x"57596871", x"430C264E",
									 -- x"716A787D", x"80799C85", x"8D814142", x"4A1A535D", x"625C6357", x"3666330F", x"30151332", x"5F3C3939",
									 -- x"3F6487BD", x"A5545568", x"7B675A6D", x"7B8B6282", x"8C9F7649", x"638FA3B1", x"1A26A992", x"7EBCA5AD",
									 -- x"979A8FA1", x"998B8C8A", x"A5A3979E", x"A4B4629F", x"B17D6462", x"565E8295", x"878B9497", x"968698AD",
									 -- x"B5B4B4A9", x"907B5C7F", x"86727D6C", x"56656467", x"6591928F", x"787A7E92", x"8FAA7A80", x"8A85A3A0",
									 -- x"A1A09B87", x"8DA6AAAC", x"AA98BD82", x"8D7A8D87", x"C6C681BE", x"7FD5A6B2", x"B1BA5D3A", x"19636B62",
									 -- x"70B7969C", x"A699B282", x"40697B79", x"4A57935A", x"4E51505E", x"5E4E6558", x"6D6C4951", x"6E636F87",
									 -- x"67546F65", x"71587A7D", x"745F514C", x"5F515060", x"605D6264", x"434F4F79", x"5F4F5327", x"6BA84F6A",
									 -- x"5A49495E", x"5F3E5B66", x"56466058", x"564498C6", x"B43E6CA9", x"535C5952", x"455F4747", x"622C4F5F",
									 -- x"54604F65", x"5E364F5E", x"5E5D7F6E", x"54485968", x"6A4D5369", x"806A698B", x"6F848B84", x"7163666B",
									 -- x"976A7C74", x"8464704E", x"4E5B5B65", x"5C505959", x"4F616870", x"685B6463", x"5C5B595B", x"58595361",
									 -- x"7C816448", x"40335D68", x"3B5B6538", x"4B696086", x"65798C6B", x"73658CA7", x"98989899", x"98999EA4",
									 -- x"ACAEAEA8", x"A29E9D9C", x"9D9B999A", x"9C9C9A97", x"9D9EA1A7", x"AAA9A8A8", x"A9A8A9AB", x"ACAAA9AB",
									 -- x"A8A5A09D", x"9DA0A09E", x"9D9F9E9E", x"A2A2A0A1", x"A4A4A5A6", x"A7A9ABAB", x"AEB0B2B3", x"B4B5B6B6",
									 -- x"B9B9B8B8", x"B7B6B6B6", x"BABDBFC0", x"C2C5C7C7", x"C6C4C3C2", x"C2C4C9CF", x"CED2D3D1", x"D1CECFD3",
									 -- x"E0E6EFF8", x"FCF8EEE6", x"EBECE9E6", x"E7EAE9E5", x"D2CFCFD0", x"CDCAC8C4", x"BAB0A39B", x"9296999B",
									 -- x"999C9E9E", x"9793928B", x"87837F7B", x"78757373", x"7274797A", x"7F838A8D", x"9EA4A3A2", x"A4A6A5A7",
									 -- x"A5A3A4A5", x"A3A6A6A0", x"9C948A83", x"7E7A7878", x"7D7C7C80", x"88979A46", x"6887695F", x"5A315477",
									 -- x"7A814465", x"775C4150", x"63444937", x"2A657564", x"6E6D6157", x"587D779A", x"7D4A4D25", x"18200012",
									 -- x"00000019", x"14212937", x"46404125", x"00092940", x"41342D2F", x"2A604401", x"21664838", x"4D494C4F",
									 -- x"4F62514E", x"4352532B", x"3F5F6444", x"5782827C", x"1D034171", x"61704E4F", x"51593B1F", x"2C6E7463",
									 -- x"64888284", x"53807C5A", x"395C425D", x"407D7079", x"856A5880", x"5342632A", x"09140832", x"5B4C838A",
									 -- x"3979796F", x"565A5F80", x"8D7BA381", x"70995E7D", x"A4AAAC8A", x"91AE9D82", x"90722868", x"AE8CA4A1",
									 -- x"98AD8095", x"9D9A8D92", x"9794A282", x"8F7D398A", x"92442C39", x"767F899D", x"98839A78", x"849A949F",
									 -- x"99ACB26F", x"6B897F75", x"6F7E7B83", x"6D7A6D42", x"3F8597A1", x"85939372", x"90969EA5", x"A1ACA69A",
									 -- x"9A8D8F95", x"9397929C", x"C19990A3", x"A8A2340B", x"958894AC", x"8B85B990", x"A9D0ADAF", x"805C7B8D",
									 -- x"6DA99DAA", x"979A9165", x"58697E6D", x"76827473", x"72696E73", x"6C73787D", x"7C7D8D95", x"78725B62",
									 -- x"63788373", x"75703C50", x"3D48463E", x"3B271B35", x"37414C57", x"5E5B5652", x"51354A39", x"4E2D6E63",
									 -- x"3E47636C", x"6A4D6959", x"715C6D70", x"7B768676", x"7B805A72", x"6A61706D", x"6D5E9099", x"605A5D5D",
									 -- x"5D5B786E", x"65545A63", x"5F56726A", x"60476A64", x"83456277", x"7A5C5E58", x"5D5F4055", x"44533B3A",
									 -- x"3D68505C", x"5961524D", x"535A5657", x"4F4D584E", x"50555F5E", x"525B6962", x"5559636B", x"655B515E",
									 -- x"7B5D3A4C", x"517D6940", x"4652414D", x"7D6E6D83", x"55748066", x"78435698", x"9A9B9C9A", x"97979DA5",
									 -- x"A9ABABA8", x"A4A29F9D", x"9B9A9A9B", x"9B9A9999", x"94979DA3", x"A5A3A3A4", x"A1A1A3A5", x"A4A09FA1",
									 -- x"9D9C9691", x"90949593", x"97979392", x"96979698", x"95969799", x"9B9E9F9E", x"A1A3A5A8", x"AAACAEAF",
									 -- x"AEAEADAD", x"AEAFB0B1", x"ACAFB1B0", x"B1B3B5B5", x"B3B3B5B8", x"BAB9BBBF", x"BAC0C0BE", x"C0C0C0C2",
									 -- x"C7C9CFD6", x"DAD7CFC8", x"CCCECDC9", x"C8CBCDCB", x"C9C3C4C4", x"BDBABAB5", x"B6AEA3A2", x"96979393",
									 -- x"939C969A", x"91868C81", x"80787578", x"77706C6D", x"676B7170", x"78798187", x"90979A99", x"9C9B9999",
									 -- x"9A9A9B98", x"95999F9F", x"968F8783", x"81808081", x"8C97999F", x"9B9FBD5E", x"1130417F", x"70276B82",
									 -- x"6C5C8A72", x"7B527965", x"56536166", x"6B7F6F82", x"97946C52", x"607C7675", x"7E777A68", x"1A000400",
									 -- x"02000913", x"163E4354", x"3C382C23", x"06002136", x"3A333F3B", x"505F471B", x"42654D40", x"373F3D2D",
									 -- x"273A4C5B", x"6B8E7A7D", x"7759606B", x"756F8062", x"2A1B1E28", x"293B5C6E", x"48211A5F", x"806B7152",
									 -- x"6E57766A", x"7657201A", x"2D8E7962", x"63878079", x"7F71597A", x"7A6C7071", x"0714151C", x"39A2977C",
									 -- x"3D51324E", x"588B959A", x"B1927A9E", x"D48B71A7", x"AFA5ACA3", x"B2A8AA9D", x"9E9D9342", x"63AE9F9D",
									 -- x"8F67463E", x"4169628D", x"B3B09189", x"8B732469", x"5A4D74A9", x"A78A9694", x"83949482", x"9592A1AE",
									 -- x"B1A9B88E", x"2C373F3F", x"6B6F6967", x"7090943D", x"279F808E", x"8C8CA18A", x"8087969B", x"96A0949C",
									 -- x"9E999D9F", x"A2A09A9A", x"A6B3A1A2", x"A3BABD58", x"84849488", x"897AA06C", x"6B627E8B", x"786C6158",
									 -- x"6D707878", x"6E797989", x"87635774", x"807C676A", x"716A896E", x"797A7895", x"6E6A6D66", x"79685758",
									 -- x"5C6A97A2", x"B3823943", x"2852474A", x"4840323A", x"53554482", x"B0267540", x"556E5574", x"646C7D61",
									 -- x"62626F60", x"6689694C", x"57646A70", x"565B5C52", x"4F355559", x"544B6062", x"6A803E3E", x"705C6269",
									 -- x"634A6157", x"5462605A", x"5E5B5864", x"2E324C5A", x"7A785E64", x"63554B3F", x"5A5F614F", x"4B3C4C4D",
									 -- x"57635C59", x"4D6D7F5C", x"594E5B59", x"4F594A46", x"525D5C4B", x"50615D65", x"63626570", x"686D6368",
									 -- x"8858537B", x"8F743C2F", x"3E535C51", x"5A6B7576", x"6A736D46", x"18276571", x"7C6E8CAE", x"9FA79DA7",
									 -- x"A8AFB1AB", x"A4A3A5A7", x"A3A2A09E", x"9C9C9D9E", x"999DA1A1", x"A1A1A09F", x"9E9F9B9A", x"9C999493",
									 -- x"99958F8C", x"8A8A8988", x"8A8B8B8B", x"8A8B8D8F", x"8E8D8D8F", x"92949493", x"92999A99", x"9DA0A0A0",
									 -- x"A5A3A3A5", x"A6A4A1A0", x"A5A5A5A7", x"A8A8ABAE", x"ACAAA9AC", x"AFB1B2B3", x"B3B3B5B7", x"B7B5B7BA",
									 -- x"BDBEC0C1", x"C1C0BDBB", x"BABABABB", x"BDBDBCBA", x"B8B6B4B2", x"B1B0AFAE", x"ABAAA8A4", x"A19D9894",
									 -- x"97949293", x"93908882", x"80777478", x"766D696B", x"686A7175", x"71747F87", x"8D939694", x"94969692",
									 -- x"97928A8D", x"8F8D9498", x"8F8A8582", x"7E7C7B7E", x"8699A5A8", x"ABABAFB8", x"96632652", x"2E637260",
									 -- x"48646F62", x"5F436F56", x"787383A1", x"6D426B7B", x"82786B50", x"7B706A65", x"54273535", x"3F000708",
									 -- x"0C0A0200", x"1E3D755E", x"23255723", x"0003002B", x"31261F1D", x"2D526403", x"8A784F5F", x"34316F88",
									 -- x"98625147", x"65555A6C", x"4C5D6261", x"84762811", x"23272321", x"1A182732", x"1A328C7C", x"6159707F",
									 -- x"85354337", x"496F6476", x"45738772", x"8461856A", x"9146537C", x"574D6320", x"31251F2E", x"43494F2E",
									 -- x"2C272834", x"39549773", x"919076B7", x"9E9FC58D", x"6995A89E", x"969FB490", x"8080B2A7", x"94789689",
									 -- x"8CA28E8C", x"823A3045", x"3E6D8089", x"8376384C", x"7CB5BEA2", x"86928D9C", x"97958E8A", x"8C8D8095",
									 -- x"9A9AABB4", x"73726251", x"2A3B5A5E", x"6D6D5D20", x"47966674", x"71768599", x"8078788A", x"8779766B",
									 -- x"7A908984", x"84879389", x"7F808682", x"8D5F7C8C", x"727D6868", x"706E7566", x"587A8A5B", x"625B5C56",
									 -- x"62626274", x"6C6D6F67", x"675B6969", x"66715E6F", x"62737064", x"74715C6D", x"626C5A5E", x"64577C83",
									 -- x"5C5A6C67", x"605C6361", x"855D5859", x"81736664", x"665C5370", x"4E4D5C64", x"60665E60", x"6D6C7089",
									 -- x"693F7B7E", x"777E8C7E", x"81645F58", x"A863655B", x"572E486C", x"81627B59", x"57837796", x"5B6B777F",
									 -- x"5F7E3853", x"6267615A", x"61616360", x"63645B5A", x"754B4661", x"5B616F74", x"446B9B71", x"6869636E",
									 -- x"60515363", x"D9FFFFC9", x"425F6650", x"4A5E5A5E", x"5F656D73", x"8895648C", x"7577747B", x"787F8E7D",
									 -- x"85707144", x"5B365153", x"41667E4C", x"64827582", x"724F0B0C", x"38867580", x"81685594", x"B8ACABAC",
									 -- x"B1B4AFAE", x"B0A8A0A4", x"A1A09E9E", x"9EA0A2A4", x"A0A1A1A0", x"9F9F9E9B", x"9C9C9997", x"98948F8E",
									 -- x"8D8D8B87", x"827F8183", x"83838382", x"82828485", x"86858586", x"88898887", x"848A8B8B", x"90949493",
									 -- x"92929294", x"95969594", x"9B99989A", x"9C9C9C9D", x"A1A0A0A2", x"A4A4A5A7", x"ABAAA9AA", x"ADAFB0B0",
									 -- x"B2B2B4B6", x"B8B9B8B6", x"B2B1AFB0", x"B2B4B5B6", x"B1B0ADAA", x"A7A5A4A3", x"A5A6A6A5", x"A4A3A29F",
									 -- x"9B999898", x"9895908C", x"877F7B7B", x"79737072", x"7B737176", x"7B808280", x"86868B91", x"918C898C",
									 -- x"8C8C878A", x"89858B8E", x"91908A89", x"8988857D", x"85919DA6", x"ADAEACAF", x"B0C4AA6A", x"476E6E5F",
									 -- x"56735A6A", x"6377367A", x"71646464", x"7089857A", x"89525566", x"60553250", x"4043461D", x"3E272743",
									 -- x"36412F1B", x"282A212D", x"12374613", x"00080421", x"472E4861", x"3C221405", x"76684540", x"2F345287",
									 -- x"6660514E", x"62525B48", x"3C434534", x"2E241425", x"1B1C191E", x"201D2221", x"16211153", x"7B5C724B",
									 -- x"056E6B75", x"9E7A6889", x"88914F5D", x"5D283329", x"40263429", x"231E192D", x"2A312734", x"3623232C",
									 -- x"291F2138", x"393F5444", x"547D8D9C", x"AC748FA2", x"859FB5B7", x"95748A9E", x"8699BFAF", x"97898A66",
									 -- x"A3A7B1BF", x"B59EA4A3", x"5D2F336C", x"AC9041B7", x"B19D8498", x"72626B85", x"84787278", x"7B887C6E",
									 -- x"6B72757D", x"9C6B717E", x"736B5857", x"736C6271", x"5661615C", x"5C646A64", x"876D6265", x"725B6B61",
									 -- x"67635454", x"595D6865", x"58645552", x"576F6169", x"5F625B5E", x"65696F70", x"786B7163", x"655E756A",
									 -- x"564A5461", x"6D686F6E", x"6868695E", x"636F6B65", x"634D5B6D", x"67676457", x"5D59555C", x"645D6351",
									 -- x"54565A61", x"7B726876", x"6E635E66", x"5F554861", x"5E5E5C53", x"5E746C8B", x"83747580", x"76716C64",
									 -- x"60566E6C", x"79757C7B", x"7B848478", x"7159616B", x"707A847C", x"7B7CA5A3", x"9D849276", x"88846572",
									 -- x"79655564", x"595E606F", x"62566063", x"5E6A654E", x"4C574E5F", x"60665764", x"6459516E", x"6F655263",
									 -- x"5C525D61", x"9C8D8F92", x"57646760", x"67737175", x"7C7C9493", x"8C8E8688", x"97978589", x"87737476",
									 -- x"3B2D3231", x"1D4B637F", x"6C93655C", x"95763C27", x"1D104885", x"967D5A69", x"4B5A5F46", x"7BAFB2AF",
									 -- x"ACAFA8A6", x"B0ADA6AB", x"A4A29F9E", x"9E9FA09F", x"9E9C9996", x"97979490", x"9495918F", x"918E8989",
									 -- x"85868582", x"7E7C7D7E", x"7D7B7A78", x"78797979", x"7E7D7B7A", x"7B7D7E7E", x"7D828282", x"878A8989",
									 -- x"82868887", x"898D8E8D", x"908C8A8C", x"8F8F8D8D", x"93929394", x"95959799", x"9B9C9DA2", x"ACB7BAB8",
									 -- x"B8B7B7B8", x"BABBB9B7", x"B1AEA9A7", x"A8ABADAE", x"ABAAA8A5", x"A2A09F9F", x"9B9EA0A0", x"A1A3A4A4",
									 -- x"A5A4A4A3", x"A2A19F9D", x"9995918E", x"8C898786", x"7E7F8383", x"7D7D8387", x"87848589", x"8A888B90",
									 -- x"8E8C8688", x"89868783", x"89939091", x"9393978D", x"91989A98", x"9BA4ADB1", x"ADAAA8CF", x"967A6772",
									 -- x"7DBC936F", x"7EBF9A77", x"9A6D7E7A", x"4F747D89", x"56624B67", x"50615D8A", x"6E615656", x"55402540",
									 -- x"404F3C48", x"54686B41", x"15010000", x"13131320", x"325A5A91", x"9197694F", x"3A1C2A48", x"4F523A4F",
									 -- x"4B575E42", x"37393C31", x"2015171C", x"1D20211A", x"23221D23", x"26211E16", x"2422140F", x"04273404",
									 -- x"46875A49", x"8277343C", x"61863638", x"301E1C16", x"27182029", x"271F2526", x"1D262028", x"202D3A36",
									 -- x"34332833", x"32261427", x"3932343D", x"6B74699B", x"73718E9D", x"7666757B", x"8291897A", x"7A7B7578",
									 -- x"645C606C", x"6969696B", x"757C4D42", x"6A5B5B68", x"4F584345", x"46263D4A", x"3F484C52", x"464A4F4E",
									 -- x"575C585C", x"7F5C656C", x"5D626A65", x"6670635E", x"6F65795F", x"5D5D6265", x"61645F62", x"635D6555",
									 -- x"635F5E60", x"5E61686B", x"69616D7C", x"6B635B61", x"70727163", x"64757572", x"6B566267", x"5A49695F",
									 -- x"595E7062", x"5D5C636C", x"716E5E52", x"58545D4F", x"5F63635E", x"575D6356", x"636E6B51", x"6466536B",
									 -- x"6D656B78", x"8B867C7F", x"6B7D9083", x"82757377", x"758D7E81", x"93847E67", x"6C849088", x"6A646A76",
									 -- x"6A716867", x"715D5C5A", x"495D5951", x"6A6C6B70", x"72758189", x"61537580", x"6D493B53", x"4B1B4A3F",
									 -- x"4B375F63", x"50626966", x"63717263", x"656F7585", x"72827A7C", x"7E8A838A", x"827F9583", x"76927A79",
									 -- x"7867807D", x"5A5F6E65", x"6F73787C", x"7B859390", x"95898387", x"929FA289", x"85959483", x"78604F61",
									 -- x"83935855", x"366C7479", x"759565A1", x"6D09585B", x"538B9087", x"698B6435", x"26616261", x"64589FB0",
									 -- x"AAB0ADA8", x"A8A9A6A4", x"A6A39E9C", x"9C9B9A98", x"9B9A9896", x"9595928D", x"8D8E8B89", x"8B898586",
									 -- x"7F7C7A7A", x"7B7A7774", x"76747170", x"7071706F", x"74737171", x"7275797B", x"7C81817E", x"81828284",
									 -- x"7F868987", x"888D8F8D", x"8D8A8889", x"8B8B8B8B", x"908F8E8F", x"8F91959A", x"9FA4A8AE", x"BBC9CECB",
									 -- x"D1D0CECE", x"CDCAC5C1", x"BAB5AFAA", x"A8A9AAAB", x"A9A9A8A6", x"A4A3A4A5", x"A2A4A6A5", x"A6A8AAAA",
									 -- x"ACACACAA", x"A9A8A8A9", x"ABACAAA7", x"A5A5A19D", x"9F9C9C97", x"8E898987", x"8A909291", x"9092908B",
									 -- x"8C8D898B", x"8D8C8E8B", x"8B938D91", x"93929A92", x"979FA29D", x"9DA4A8A4", x"ACB1B7BE", x"756D7F6C",
									 -- x"72827991", x"80747B4A", x"80B79D87", x"66693C2F", x"2A66626B", x"84724E2B", x"5A191B5B", x"373A3316",
									 -- x"39434B5B", x"6682723B", x"273F160F", x"0E0B427D", x"33825276", x"9B913932", x"3115262F", x"23261E23",
									 -- x"19182518", x"16292520", x"151E272A", x"1D223328", x"30312E33", x"3431322E", x"30333439", x"251F1925",
									 -- x"26271525", x"4950321C", x"55663E25", x"231F192B", x"2C261E1A", x"12323528", x"2829323F", x"2D2B3530",
									 -- x"3739383A", x"34332C3F", x"343A484B", x"5A584D5F", x"4F575E5B", x"5664584F", x"5D53555F", x"57565554",
									 -- x"54534A4B", x"494F4844", x"3343554E", x"4C544E45", x"4037353A", x"38224336", x"414A3B47", x"5049444C",
									 -- x"4D4A585A", x"52545453", x"614C6258", x"3E536765", x"52535450", x"50525B5A", x"555F605A", x"535D5951",
									 -- x"59616A5F", x"53534D45", x"586A7169", x"6F4C6169", x"5D728275", x"686B6A68", x"71646A69", x"67697869",
									 -- x"565E6C62", x"58655966", x"6D747377", x"817D806F", x"508B8D81", x"8D897971", x"70867F8D", x"8F808B79",
									 -- x"87808B8B", x"82838178", x"7686827F", x"8494867D", x"7B796767", x"6C5A615C", x"5F6B605F", x"61655D67",
									 -- x"68635864", x"64596057", x"6A847072", x"7D7D7D93", x"73718799", x"8790886C", x"78777778", x"777C7B7C",
									 -- x"637E836D", x"7B888488", x"8E818584", x"7F868A8A", x"898E9B9A", x"A19BA1A2", x"92A0A2A2", x"A0917F95",
									 -- x"95998F85", x"9BA691A5", x"A3B19696", x"A2A69792", x"8F8C7A7F", x"7A868F8C", x"686D7E5E", x"5C71595C",
									 -- x"4138597B", x"6671686D", x"73697D73", x"6D6CA591", x"73848499", x"7A7C6358", x"656F7471", x"64656CB0",
									 -- x"B8B5BBBD", x"B6B4B4AB", x"ABA8A5A4", x"A5A6A4A3", x"A0A1A19F", x"9D9A9692", x"8A8B8783", x"83807D7E",
									 -- x"7D7B7878", x"7A797471", x"6D6B6A6A", x"6B6B6B6A", x"6B6D6F71", x"73767A7C", x"7F848482", x"8283868B",
									 -- x"8A929795", x"94979895", x"9F9D9B9B", x"9A999B9E", x"9B989696", x"989BA2A9", x"B2B7BCBE", x"C5CED0CC",
									 -- x"D4D4D4D4", x"D2CDC6C0", x"BFBBB5B1", x"B0B0B0B0", x"AEAEADAC", x"AAA9A9AA", x"AAABABA9", x"A8A9A9A9",
									 -- x"A8A9AAA8", x"A6A5A7A9", x"AFB2B2AF", x"AEB0AFAA", x"ACAAAAA6", x"9E9D9F9E", x"9B9FA09E", x"9EA1A09B",
									 -- x"93989695", x"908A8D8D", x"8E8D868C", x"91909590", x"92949699", x"9A938C8B", x"84838E88", x"73796560",
									 -- x"696E8858", x"72949482", x"72667950", x"1D302450", x"717B7F6A", x"606E4D67", x"53225F69", x"52597D28",
									 -- x"35606974", x"5F795D0A", x"2846133E", x"34458284", x"57515E53", x"4820070D", x"0C1C2326", x"27283022",
									 -- x"2B2E242B", x"282C392F", x"35383135", x"3A425046", x"42464346", x"47454642", x"3A463A41", x"3F393C3A",
									 -- x"301A1F22", x"22202937", x"4B372F1C", x"2B261623", x"203A3727", x"75E04729", x"3E3F3325", x"28222628",
									 -- x"251B323C", x"3A445043", x"8895524A", x"5348565A", x"51495B59", x"3F53584F", x"51565149", x"4F504E4F",
									 -- x"424D4D54", x"4B585B41", x"3660423E", x"32514433", x"43383954", x"3B384146", x"504D3648", x"5D59463F",
									 -- x"45384C58", x"59393B54", x"3A3B4E30", x"2A384442", x"44494E58", x"4B4E5C4C", x"523E4B3C", x"4E4C484D",
									 -- x"51565B59", x"616E675A", x"5A5A5D63", x"605E7868", x"6D635864", x"73747472", x"6B626D54", x"45637E81",
									 -- x"493C474A", x"4B5E628B", x"7A868275", x"72848175", x"5A736B6A", x"77736F6E", x"6D606567", x"5E64655C",
									 -- x"61686F67", x"5D606063", x"5D5A515B", x"6D71645C", x"57675B54", x"5859565F", x"5F585661", x"5E5C5D69",
									 -- x"6E5B5360", x"5C5A605E", x"66636A6B", x"88616F57", x"5C647B77", x"77897B88", x"8C908A85", x"95A1A5A7",
									 -- x"B8B19D8F", x"8B8B90A0", x"96858D97", x"9089878B", x"8388887E", x"84777E8E", x"80756A80", x"68716E82",
									 -- x"716E7859", x"616D7475", x"747F7584", x"74838885", x"9096A9AF", x"8D8BA5BF", x"B9ABB69A", x"87A19F92",
									 -- x"3E3F2325", x"262A4755", x"547B7363", x"928D122B", x"8A90979D", x"646D6B86", x"66996E47", x"738C45B8",
									 -- x"D3C5C8D2", x"CECCCECB", x"C0BFBEBE", x"BFBFBEBC", x"B2B3B3B1", x"AEABA7A3", x"9C9C9690", x"8D888384",
									 -- x"7B7C7C7B", x"78757372", x"70707071", x"73747474", x"74798084", x"8687898B", x"92979897", x"999B9EA4",
									 -- x"A7ADB1B1", x"AFB0AFAD", x"ACAAA8A7", x"A5A3A5A8", x"A9A6A4A4", x"A5A9AFB5", x"B2B6B9B9", x"BCC0C0BE",
									 -- x"C4C6C8CA", x"C9C5C0BC", x"B9B7B5B4", x"B5B6B6B5", x"B5B4B2B1", x"AFADABA9", x"A7A7A5A2", x"A1A1A09E",
									 -- x"A1A2A3A2", x"A0A0A1A3", x"A9ABABA7", x"A8ADAFAD", x"A9A9AAA5", x"9C9B9FA0", x"A6A3A3A5", x"A2989190",
									 -- x"96938E93", x"948D8C88", x"88878888", x"85828387", x"8A8C8C8D", x"856E6A7E", x"70655A64", x"777A6B7D",
									 -- x"7A714457", x"66554059", x"71474546", x"5C6B8A79", x"6B6C726F", x"677A3C58", x"6F525C43", x"35526A3C",
									 -- x"274E4539", x"669B2C21", x"261E0514", x"37302D3E", x"28180517", x"254C5A6E", x"88683A2D", x"2F2B4732",
									 -- x"27303230", x"2A2F3B3E", x"3E3F3539", x"3C333435", x"33353338", x"3D3C3A32", x"3A3A4645", x"4046483F",
									 -- x"3F3D303A", x"371C3A40", x"39352F25", x"2624150A", x"16364442", x"8B733A3D", x"34332E1B", x"242B2914",
									 -- x"1C1A2E30", x"51544F46", x"866F292E", x"4F605253", x"44495151", x"50514A56", x"58536766", x"5D5F6952",
									 -- x"5F655C63", x"5C4E4B45", x"3444452C", x"364B3034", x"272F3742", x"312B1B2D", x"3A404652", x"4D4F493C",
									 -- x"2948514F", x"5E5D6E60", x"5B525C52", x"5E51515D", x"52586158", x"58535659", x"5549574C", x"5C635961",
									 -- x"6A675E60", x"69675F5A", x"5E59606A", x"796B6376", x"626B6B77", x"7F736D6E", x"74494C37", x"20444F44",
									 -- x"32212E20", x"20283656", x"3E4B5957", x"4F5A4947", x"5B5E575A", x"60574F4E", x"53544D58", x"5856554E",
									 -- x"413F4A50", x"4853595A", x"565A5F58", x"644B4942", x"46423D4F", x"515E5757", x"60625D58", x"5E5D5C60",
									 -- x"6D656064", x"6860555E", x"606E6066", x"67606666", x"658B656E", x"70666D2D", x"3268694E", x"4F504439",
									 -- x"51607867", x"5A827861", x"7567616C", x"7D76656C", x"65696C7A", x"737C7B7C", x"7E788B7A", x"6E969584",
									 -- x"758BA390", x"72786E5C", x"6969696C", x"393D566A", x"6D555456", x"6E63595C", x"6F677177", x"5849574B",
									 -- x"472F3336", x"37262826", x"3C3D314B", x"756B9141", x"307BAC67", x"6053603F", x"46586868", x"6D584D94",
									 -- x"D6D7D4D2", x"D5D4D2D5", x"D4D4D4D3", x"D2CFCDCB", x"C7C6C4C3", x"C3C3C1BD", x"BAB9B2AB", x"A7A19D9D",
									 -- x"9C9D9E9D", x"9B999796", x"8C8D8F91", x"91919192", x"94989EA1", x"A1A2A4A6", x"AEB1B2B4", x"B8B8B8BB",
									 -- x"C0C2C5C6", x"C5C4C2C2", x"C3C1BFBF", x"BEBCBCBD", x"B8B5B3B4", x"B5B6B8BA", x"B0AFAEAE", x"AFB1B2B2",
									 -- x"B9BCBFC1", x"C0BEBBBA", x"B2B1B0B1", x"B2B3B2B1", x"B3B1AFAE", x"AEABA7A3", x"A4A2A09D", x"9D9D9A97",
									 -- x"999B9C9C", x"9B9B9C9E", x"A2A4A3A1", x"A3A8ACAC", x"ABA7A6A8", x"A8A9A398", x"8E7D6A5E", x"57576069",
									 -- x"746D6671", x"78767A7B", x"87838B85", x"858B868C", x"828F887A", x"7466657C", x"77787558", x"61405D6E",
									 -- x"63445E71", x"85716AA1", x"827F9889", x"9677786F", x"656E6A59", x"766A6B5D", x"475E817D", x"84477472",
									 -- x"5B441A1E", x"434C1224", x"12276C61", x"784E0605", x"113C7C94", x"B092A99A", x"76523832", x"35273D37",
									 -- x"34334138", x"3E443333", x"3B383239", x"413E3B3D", x"31343136", x"3D424640", x"455B3D3A", x"4A413B36",
									 -- x"3A384C44", x"2F222237", x"393D3137", x"32333337", x"3C3E4543", x"365D4247", x"331A1B1D", x"0F0D1718",
									 -- x"07162D15", x"3C422F3E", x"201C4541", x"59575565", x"514C5457", x"5C5C564B", x"5555595A", x"5C535050",
									 -- x"4B4A474B", x"55484655", x"604C654A", x"4933202C", x"3D223543", x"39383F41", x"3C404A51", x"4B524B45",
									 -- x"4A4B4960", x"5C566460", x"5B5C6154", x"575C6154", x"514F4B40", x"58534E5C", x"666D665C", x"5E6F696A",
									 -- x"747C7682", x"8D838795", x"8D848976", x"72626263", x"5E686259", x"66655354", x"472B3537", x"22363E40",
									 -- x"392E3F3C", x"4854514B", x"4E4C5A5A", x"53514955", x"4F595850", x"52524A4F", x"53434D59", x"4F626251",
									 -- x"544E5358", x"51615B4D", x"3A534C55", x"464E5161", x"39425442", x"3F79684B", x"454D4F40", x"47444745",
									 -- x"3946494C", x"5A524C55", x"3F55584D", x"605E565F", x"68545A62", x"59676065", x"5B545B74", x"615C6C5D",
									 -- x"5B575449", x"585E466B", x"655A6767", x"585B6059", x"625B5B6A", x"52636A6B", x"61583C26", x"4E425A60",
									 -- x"6B6A636A", x"686B646A", x"70756660", x"686A6A89", x"6E737369", x"85757084", x"6F6F7A91", x"94847D7B",
									 -- x"50614C54", x"43484449", x"36392C47", x"28327232", x"43416984", x"7F5D9071", x"383F6357", x"6C415C4A",
									 -- x"AED0D3C7", x"D2D6CED0", x"D4D5D6D5", x"D2CFCCCB", x"C8C5C2C2", x"C6CBCBC7", x"C1C1BBB4", x"B1ABA7A9",
									 -- x"B3B1AFB1", x"B5B6B2AD", x"ABAEB0B1", x"B0AFAEAF", x"B0B2B4B4", x"B3B5B9BD", x"BEBFBFC1", x"C7C6C1C1",
									 -- x"C5C5C6C8", x"C8C6C5C5", x"C7C4C3C4", x"C6C4C2C1", x"C3C1BFC1", x"C1BFBDBD", x"BFB9B2AF", x"ADACACAE",
									 -- x"AEB0B2B2", x"AFAEAEAF", x"B0AFAEAD", x"ADACAAA8", x"A9A7A6A7", x"A8A7A29D", x"9F9D9997", x"9898948F",
									 -- x"94959798", x"97989899", x"9D9FA0A1", x"A3A6A9AA", x"A4A8A899", x"7D655347", x"4D535758", x"5D62625D",
									 -- x"52504C4D", x"443B4958", x"55475054", x"70908684", x"858D6B48", x"566C7582", x"6F6D6C66", x"797B585E",
									 -- x"6C787D7D", x"6A758386", x"87808764", x"726A6791", x"606A6B8A", x"7467856A", x"68844B87", x"694D90A1",
									 -- x"BBA88849", x"29112636", x"317BA1A8", x"A9752537", x"34474123", x"1921101A", x"1E2B2C1E", x"423E3C4B",
									 -- x"41463E3A", x"3F343B3C", x"3B3E4244", x"494C4740", x"49493F3B", x"3A3D4748", x"473F293E", x"48413835",
									 -- x"343A2F3A", x"322A2C33", x"3640383A", x"48594941", x"454A4545", x"3C444436", x"342C242F", x"38413637",
									 -- x"3C47794C", x"43564E58", x"5E67605D", x"4F443E44", x"3B3E3D3A", x"49444446", x"48474649", x"48464342",
									 -- x"453C5041", x"3B494C3C", x"4B4B3D4E", x"4D404041", x"49575551", x"3D48464F", x"5D574F53", x"5F624E5B",
									 -- x"635D635E", x"65676A6E", x"6A6B696D", x"69616265", x"6B67676F", x"63596870", x"75776F6D", x"857C7F71",
									 -- x"74827072", x"76626776", x"59604648", x"5550514B", x"4C4D4E44", x"56594053", x"66594E53", x"4A494250",
									 -- x"66545356", x"4C595558", x"54565E52", x"4F4A4D50", x"473F4339", x"333D3F43", x"5A7F6666", x"50405654",
									 -- x"56695542", x"4B512D20", x"28373341", x"3830364A", x"56613942", x"371D3548", x"34153248", x"4A425445",
									 -- x"3D4D4F4C", x"504A5554", x"42475A50", x"454E3639", x"4451585C", x"525C5376", x"673A3A4D", x"62535B5F",
									 -- x"64515B66", x"6A63565D", x"6861523D", x"42596061", x"4A606F79", x"71687092", x"64535F42", x"38425647",
									 -- x"4F616C4A", x"644F6264", x"6D55635F", x"5E646148", x"62666567", x"69686862", x"61686E5B", x"696B4D64",
									 -- x"4F5D5E5D", x"41434943", x"574E594F", x"2436643C", x"41505B65", x"585C76A0", x"6C666480", x"6D48665E",
									 -- x"8CCBC5C2", x"C5C7C6CB", x"C9CCCAC9", x"CDCDC7C4", x"C4C4C1BF", x"C0C3C5C5", x"BBBDBCB3", x"A8A2A3A7",
									 -- x"ADAEB1B5", x"B7B6B1AD", x"ACB1B5B6", x"B6B5B3B0", x"BABEC3C6", x"C7C9CCCF", x"CBC8C9CD", x"CCC7C3C3",
									 -- x"C5C5C5C5", x"C5C6C6C6", x"C5C6C3BF", x"C1C5C5C2", x"C5C0C0C4", x"C3BFC4CE", x"D6CCC2BA", x"B3ADADB1",
									 -- x"ADAAA8A8", x"A9A7A29E", x"A2A19F9F", x"A0A1A2A2", x"A09F9D9B", x"9A9A9DA1", x"99979094", x"968F9196",
									 -- x"97929592", x"97909494", x"9895A39B", x"97A29EA2", x"9EAE9038", x"3B4A333D", x"45424642", x"4D4A5548",
									 -- x"3C4D424D", x"45514A40", x"1812141A", x"045C968A", x"8C8B7937", x"2C303E4B", x"64836C71", x"7E605D5F",
									 -- x"6C745774", x"7A7E507C", x"947D905F", x"6E735E84", x"6C496980", x"4E6C7377", x"756B5F5E", x"7D8A729C",
									 -- x"998AA09C", x"8E7E64A5", x"59241021", x"251F534B", x"2E213030", x"2F34282E", x"2533322F", x"4639403E",
									 -- x"3A403C46", x"3E383C3F", x"43494B41", x"45424543", x"4B3C383C", x"3D38363B", x"2E3F3439", x"3E404246",
									 -- x"40484133", x"39473C42", x"42474746", x"4848484F", x"51505263", x"594F4B4C", x"49525C50", x"65656A4F",
									 -- x"494D524D", x"4E524E50", x"51526059", x"5259544F", x"564F5151", x"494F5753", x"58595250", x"4453505F",
									 -- x"646F6281", x"796C6077", x"705D5A69", x"61776B71", x"6B5D695C", x"82AFA379", x"90CA9577", x"786F6A60",
									 -- x"6E6C716A", x"6A747D72", x"707C6C77", x"7D788A75", x"7A908781", x"838F9165", x"6A70695E", x"6E5D615A",
									 -- x"66645F5A", x"5C595654", x"52555659", x"50585754", x"56618E55", x"606B6458", x"695E5E58", x"606A615F",
									 -- x"5A606455", x"5A5C595E", x"6575815F", x"56544A44", x"4F4E4B46", x"574D4044", x"4D544F58", x"4E4B4F59",
									 -- x"56535642", x"59514557", x"624D4348", x"33111221", x"3D3B1522", x"3F4E2D3F", x"3C304051", x"55585451",
									 -- x"394B3D47", x"453A444E", x"4B5E6156", x"5751585A", x"614D6867", x"645E4D7B", x"5D4C5E50", x"61554E4B",
									 -- x"65535D61", x"4D58735E", x"675F585F", x"4A645E68", x"6D6E7A78", x"7B6B6269", x"6A738B82", x"8E8871AA",
									 -- x"778D8E8D", x"93706965", x"5F6B597E", x"6A707558", x"5F62626A", x"7767664C", x"5C68645E", x"707B4150",
									 -- x"5041677F", x"5D636348", x"584D445D", x"442A3B4C", x"4842123A", x"6A35565F", x"7894647A", x"875E5B80",
									 -- x"4BA9CFB8", x"C2BDBDC2", x"BEBFBCBA", x"BEC0BEBE", x"BEBEBCBA", x"BBBDBDBC", x"B9BAB9B5", x"B1AEAFB1",
									 -- x"B1B1B2B4", x"B4B3B1AE", x"AEB0B2B3", x"B7BABBB9", x"C3C5C6C6", x"C5C5C7C9", x"C9C6C7CA", x"CAC5C3C4",
									 -- x"C5C4C3C3", x"C3C4C5C7", x"C2C5C7C6", x"C4C4C2C0", x"C4C3C4C5", x"C2C1CCD9", x"DEDCD3C3", x"B4ACACAE",
									 -- x"B5ADA7A5", x"A5A39F9D", x"98999B9C", x"9C9A9794", x"99959190", x"92939392", x"8F918F93", x"93948E8F",
									 -- x"908F958F", x"8E8F9096", x"9691979B", x"9A9A9898", x"9C995450", x"43444544", x"493D4144", x"402D3738",
									 -- x"51495447", x"3D463220", x"0F081610", x"041DA27E", x"888A8D4E", x"35354C77", x"83673A3F", x"283A5E5C",
									 -- x"66556C70", x"8387808F", x"73747D6A", x"58656070", x"66566F72", x"4D524D4B", x"5743484E", x"61635059",
									 -- x"4A484938", x"2F3A2328", x"2C213731", x"32291E22", x"34292F2B", x"2A33333E", x"43394A48", x"3E363E36",
									 -- x"3219443B", x"3F47414D", x"4647404F", x"494A3D44", x"3C40502A", x"414F4B4E", x"554E5153", x"434D524D",
									 -- x"4D454449", x"4E4E4A48", x"48574B44", x"4F4C4954", x"524D5056", x"5C565A43", x"4F4A5B57", x"3C395C53",
									 -- x"43323F60", x"6A415767", x"5C5C4A4B", x"5B616566", x"64697172", x"6A6B7171", x"858E7887", x"81756861",
									 -- x"7E7A896E", x"7077656A", x"62625960", x"58525750", x"567B85A9", x"B4999C77", x"5E647CAE", x"A6594558",
									 -- x"656C5846", x"4D575741", x"46344C53", x"45514845", x"4257443B", x"483E454B", x"44585B40", x"4C565850",
									 -- x"4C52605B", x"60545857", x"5D645E58", x"575B5654", x"53555B5D", x"50613B36", x"42565253", x"5F57625D",
									 -- x"5A655E4F", x"634F4A59", x"798CA990", x"4A6A5F64", x"65625669", x"65526350", x"594E4B57", x"5053524E",
									 -- x"60606256", x"645B5B5B", x"655F585B", x"59545754", x"56614F53", x"585F5E52", x"5A615F60", x"5D5F6757",
									 -- x"565A5957", x"6D5A4068", x"58585F5C", x"5A607162", x"5554737C", x"6E635E53", x"5D887666", x"7287687A",
									 -- x"8A8E728F", x"AE674B55", x"6555505F", x"606B8168", x"7A858474", x"54658289", x"7F5D656C", x"817D7477",
									 -- x"6F615059", x"6C817564", x"655B5C6C", x"686D7A6D", x"6F777E7C", x"63547D6D", x"5A5C6469", x"5B615F71",
									 -- x"6A666864", x"40578881", x"52675E36", x"32345A77", x"99933B21", x"1B3F5652", x"6DAEA67F", x"672C5E6A",
									 -- x"487EBCB9", x"BDBEB9B9", x"B9BAB7B4", x"B8BABABC", x"BABABAB9", x"BABBBAB7", x"B8B6B5B6", x"B8B9B8B7",
									 -- x"B6B5B4B3", x"B3B2B3B3", x"B1B0AFB1", x"B6BDC0C0", x"C5C5C5C4", x"C3C2C1C0", x"C1BFBFC1", x"C1BDBCBE",
									 -- x"C0BFBEBD", x"BDBFC2C5", x"C5C6C7C6", x"C3C1C5CA", x"CDCDCBC9", x"C7CBD7E2", x"E3E5DFD0", x"C3BDB8B4",
									 -- x"B4B0ACAA", x"A2999496", x"8F8F8E8F", x"90909090", x"8C8C8D8B", x"8A888786", x"87858682", x"808A8286",
									 -- x"8A898B8A", x"8A928784", x"8C8F8E94", x"93939B97", x"88724C3A", x"505D385C", x"5E473B3B", x"38394A4B",
									 -- x"404E4350", x"48330D0C", x"080F0414", x"02498581", x"84808573", x"6D79907C", x"57212629", x"22263F80",
									 -- x"82827787", x"653C676F", x"6C595E6B", x"5763696D", x"69595039", x"34363C3C", x"47363933", x"362B282C",
									 -- x"3128242A", x"272E302E", x"2E2E3026", x"2E322A30", x"33373836", x"3E4A4230", x"3E2C3435", x"393B3335",
									 -- x"4543404B", x"414F4B45", x"443F3B3A", x"3D363335", x"2A1E2423", x"35313C2B", x"2F2D2F22", x"13201E25",
									 -- x"2D42333B", x"2D4F5057", x"504E4D5A", x"59556161", x"5C756A73", x"6E615E65", x"6969596B", x"7C695E56",
									 -- x"7570756B", x"647D7D7D", x"71807E75", x"7A878B83", x"97948C88", x"8A8A8681", x"7D716762", x"606A586C",
									 -- x"5E584C64", x"5C455C51", x"5B5E515C", x"4D4C4C73", x"AA8D4D5C", x"37343233", x"42245B6A", x"82797FB8",
									 -- x"9A99AFA4", x"A097A08D", x"7E6A6149", x"494C3E4C", x"4746424D", x"5646515D", x"555B5D49", x"4C57535B",
									 -- x"55565F6D", x"414F5859", x"4854534C", x"56575558", x"5E4B3B51", x"4D565469", x"635A6661", x"52636863",
									 -- x"63616458", x"5C626563", x"5A514765", x"60616455", x"5C5E736D", x"574F4C6A", x"6C5C6368", x"565B6261",
									 -- x"595F635A", x"5A53625C", x"5F625F5F", x"5B596267", x"98665D65", x"6360625A", x"63706971", x"6C5E6457",
									 -- x"61606160", x"576A6152", x"5758534D", x"55535751", x"4C4B4E55", x"5F55616D", x"69656769", x"6D63636B",
									 -- x"626468A1", x"63547181", x"6E556550", x"52676948", x"56544D5C", x"5A69715D", x"7A675864", x"653D4169",
									 -- x"5F555F52", x"5A5A595B", x"62638062", x"5A63596D", x"7E7E6F6F", x"765D7389", x"7D64616C", x"675C7678",
									 -- x"49497571", x"4B3E4B69", x"6072956A", x"6699461F", x"2335405C", x"69463D38", x"28505E62", x"51425277",
									 -- x"5245ACC9", x"BBB7C2B7", x"BABDBBBA", x"BCBBB9BA", x"BABBBBBB", x"BBBCBBB9", x"B9B6B5B6", x"B9BAB8B6",
									 -- x"B7B6B5B3", x"B2B3B5B6", x"B5B4B2B2", x"B6BCBFBF", x"BCBDBFC2", x"C3C2BEBB", x"BAB9B9BA", x"B8B5B3B4",
									 -- x"B7B7B7B6", x"B6B8BCBF", x"C3C2C3C5", x"C3C2C9D2", x"D9D8D3CF", x"D2DAE1E4", x"E9E7E4E3", x"E3E0D6CC",
									 -- x"C3BBB5B3", x"ADA29C9D", x"96918B88", x"88898988", x"8A898989", x"8A8A8885", x"837F9089", x"878B8489",
									 -- x"808A8687", x"81898A89", x"898E8E8A", x"8E989380", x"6955453B", x"41453D47", x"4837313E", x"3F45504B",
									 -- x"535D5948", x"3A090B0B", x"0D140A07", x"14846F7F", x"74727E6D", x"81835B49", x"2023281A", x"517F697B",
									 -- x"7B747B6B", x"526B5270", x"825D734C", x"5E617457", x"3A3A3932", x"413C3F39", x"343B3937", x"3E323441",
									 -- x"413E3F3E", x"3C363E3B", x"3E3F3D3C", x"35374245", x"4F392430", x"392D2A2A", x"272E3538", x"3F3F3B4B",
									 -- x"3E3A3B3E", x"463E3423", x"392D2822", x"30282826", x"33282933", x"2A2E2625", x"2E282D3C", x"3B3A3546",
									 -- x"4A384B4C", x"3E3E4838", x"565B564D", x"43597157", x"4D595360", x"4F495756", x"4E4F5958", x"6F3D4A45",
									 -- x"44475C5A", x"44594F74", x"705B6C64", x"667F6035", x"5E5A4C4B", x"5D66605D", x"69665960", x"5A5E6262",
									 -- x"5E545C4B", x"48585A74", x"6D757DA9", x"92899893", x"907A6970", x"84766A76", x"5E98A66F", x"93A1AB8F",
									 -- x"9D9EACAC", x"809293AD", x"B1B0A0A7", x"7B7A6848", x"4F474951", x"4A4E5245", x"57535156", x"5758505E",
									 -- x"5A5C5D5D", x"5F5B5757", x"5C5F6259", x"5B525355", x"5A65625E", x"605A6457", x"54515469", x"56686F68",
									 -- x"63635D5A", x"6273686C", x"64626259", x"66616C73", x"65707467", x"6E8C7D76", x"7262686D", x"64676763",
									 -- x"696B7069", x"6A677477", x"69655C5F", x"635D5851", x"545A5661", x"4E405D4E", x"42575B4F", x"52626459",
									 -- x"535C614E", x"455D5D44", x"4A4F515F", x"786B5D54", x"5D5E5F5D", x"745D4B66", x"6D5B5E5E", x"56525A45",
									 -- x"44554444", x"485D616A", x"6262605B", x"4D395365", x"656E6551", x"5F655F46", x"47564B56", x"576D6145",
									 -- x"5F626061", x"5F664C49", x"626A665E", x"72755C6E", x"6B6B5C6E", x"A1825A6D", x"8890665C", x"5B73715A",
									 -- x"523A4B5B", x"75697658", x"65526257", x"615A4E49", x"3230538D", x"59777D7D", x"5441264D", x"7C666239",
									 -- x"2258CAB7", x"C0BBBEBA", x"BABDBCBC", x"BEBBB7B9", x"BBBCBBBA", x"BBBCBCBA", x"BBBAB9BA", x"BBBAB9B7",
									 -- x"BAB9B8B7", x"B6B6B7B8", x"B8B9B9B8", x"B8BBBDBD", x"B9BABDC1", x"C3C3BFBC", x"BABABBBB", x"B8B5B3B3",
									 -- x"B2B4B4B4", x"B4B4B6B8", x"B9B7BCC3", x"C5C4C8CF", x"DADCDAD7", x"DBE3E8E7", x"EAE4E2E9", x"F0EDE4DC",
									 -- x"D4C3B4B1", x"B2AEA9A6", x"A6A29E9E", x"A0A19F9C", x"969C9F9D", x"99989797", x"9A7F7E5F", x"58586678",
									 -- x"80866B66", x"5D636F69", x"7A77807D", x"8894795D", x"49391B3F", x"443D413A", x"40394257", x"4E404C59",
									 -- x"594E5C41", x"00101D13", x"11141400", x"32857D7D", x"71676B7F", x"6F362116", x"20473564", x"6F796967",
									 -- x"736C6375", x"81786670", x"6E564B4B", x"363A3235", x"363A3D3F", x"3F384345", x"444C4044", x"46444248",
									 -- x"3C39433D", x"4A434041", x"463C433B", x"38433E42", x"434A3B3A", x"403F4036", x"39342D34", x"36332D1C",
									 -- x"222E2E30", x"42413D32", x"3F433D43", x"38362F3B", x"3A304B45", x"394C36A2", x"EB823845", x"46413F35",
									 -- x"473F483F", x"4A49414B", x"40413639", x"3E383E45", x"444B4542", x"6951554E", x"49412D4E", x"38231823",
									 -- x"112D3D3E", x"4B4F5663", x"58415552", x"46565655", x"44504D4B", x"55575357", x"564E4C56", x"4F5A5F48",
									 -- x"504E6F7B", x"828CBBB0", x"9AACCAA2", x"B5A49092", x"91549492", x"9BB7A2BE", x"B1B69472", x"A79B8E6E",
									 -- x"808F9284", x"9891868B", x"9A96A47C", x"443E4D50", x"67584E55", x"494F494D", x"4B55505A", x"56575350",
									 -- x"524C5B5B", x"5D5B6B6A", x"5D525E64", x"61555850", x"58635967", x"696A7066", x"5B646A6D", x"706C5272",
									 -- x"7D69596A", x"73676D63", x"66726D77", x"7C877865", x"75666A6E", x"58616F78", x"6A676D6F", x"6A605959",
									 -- x"65626B67", x"72726B78", x"74756762", x"6B706E65", x"65625E67", x"6B776A70", x"725B6B6D", x"7A82656F",
									 -- x"6E597B5E", x"63635866", x"6460666A", x"6A64634C", x"636C6559", x"72746668", x"51656351", x"675E5B57",
									 -- x"5C61686C", x"66716942", x"5572635B", x"7670757A", x"7F7E948E", x"89706376", x"70716B85", x"92A08E8F",
									 -- x"74768E76", x"77708676", x"7CA37A6C", x"83929964", x"5F747686", x"8875665E", x"71786E69", x"7C6F6563",
									 -- x"535C4D4D", x"42765055", x"6D93685B", x"525F7768", x"6345418A", x"47624874", x"5775483F", x"7F7C9A89",
									 -- x"548ACCC1", x"BEC2B5BF", x"BDBEBCBC", x"BFBDBABD", x"BEBEBDBC", x"BCBEBDBC", x"BEBFBFC0", x"BFBFBFC0",
									 -- x"C2C1C0BF", x"BEBDBDBD", x"BCBEBFBE", x"BDBEBFBE", x"C0BFBFC1", x"C2C3C2C0", x"BCBDBFBE", x"BBB8B6B6",
									 -- x"B3B6B9B9", x"B8B7B7B8", x"B7B4B6BC", x"C0C2C6CC", x"D0D8DEDC", x"DCE2E9ED", x"ECE6E3E7", x"E8E3DFDE",
									 -- x"D0C8BEB8", x"B4B0ACAA", x"A9A6A4A3", x"A4A5A4A3", x"B0AAA4A5", x"AAA5917C", x"6144412E", x"2E354E5F",
									 -- x"585D453B", x"2F2F3F3B", x"4C485D61", x"6974625B", x"60585958", x"54413346", x"43464C4F", x"483F5364",
									 -- x"46503106", x"18150C17", x"13110B00", x"58826F6E", x"6D7C6632", x"37536589", x"8690687B", x"6C5D5958",
									 -- x"53625A5C", x"5447472E", x"2F3F3D37", x"3F3E4C3E", x"423F454F", x"463E4242", x"4444424A", x"3E474E4A",
									 -- x"4944493F", x"43423A45", x"4A494039", x"47493D35", x"3137313D", x"4C474441", x"4249413F", x"423D453F",
									 -- x"3F373D62", x"504B5151", x"4754534D", x"53616058", x"4C694248", x"50494D42", x"45261438", x"44434743",
									 -- x"3F4C3942", x"4760383D", x"3F47453F", x"45484549", x"57475156", x"50354B5C", x"48261F2A", x"2B020006",
									 -- x"211F1D29", x"444B3F47", x"575B5056", x"584F514D", x"4E5E5E55", x"534E4A50", x"312B4A50", x"495A4E38",
									 -- x"339AB69E", x"9C938799", x"9DA09879", x"A9A3A08C", x"956E87B7", x"90968B86", x"97A3BB97", x"989B7E71",
									 -- x"6A806971", x"6B5F6C77", x"6F7D634B", x"3E2A4657", x"9B9AB4CB", x"B9B58B65", x"676F6369", x"61636966",
									 -- x"616F6762", x"63626682", x"83656369", x"69738888", x"95948F9C", x"93827A78", x"8D98757D", x"947D99B5",
									 -- x"A0A77873", x"AB878E90", x"8FAF8A8F", x"8C867E78", x"697C8B85", x"7B88867C", x"7781878B", x"8D8594A0",
									 -- x"6E71827D", x"7D74647A", x"747D7A7E", x"827A797D", x"6F8C737D", x"7B887469", x"77749988", x"7A7C5D6A",
									 -- x"7A717068", x"6379646E", x"8C5E516F", x"7D616473", x"7C967975", x"969E9891", x"757A9598", x"957F8386",
									 -- x"84958DA2", x"888C9D81", x"8C9C957A", x"907B6F88", x"7F758E92", x"82938E9B", x"979C8C79", x"93968B9E",
									 -- x"8D798C9D", x"7F8A9E8C", x"8A879493", x"9492AB94", x"98A38398", x"7E7A8D73", x"746D726F", x"8379726C",
									 -- x"4B575943", x"5B443B47", x"474C523E", x"49515A70", x"615B594C", x"5C668957", x"3A407E4C", x"74497C9E",
									 -- x"B17F96C5", x"BCBBBEC3", x"C0C0BEBF", x"C3C1BEC0", x"BFC0C0BF", x"C1C3C3C2", x"C2C3C4C4", x"C4C4C5C6",
									 -- x"C7C5C4C4", x"C4C4C2C0", x"BFC1C1C0", x"C1C3C3C1", x"C3C3C2C2", x"C2C2C2C2", x"BFC1C1BF", x"BCB9B8B8",
									 -- x"B6BABEC0", x"BFBEBFC0", x"C1BDBABA", x"BCBFC5CB", x"CBD4DBDB", x"DBDFE6EB", x"F0EEEBE9", x"E6E1DFDE",
									 -- x"D0D2D2D0", x"CDCAC4C0", x"C7C7C4BC", x"B3ACAAAA", x"A3AAA794", x"7D6E6969", x"553E312F", x"30425357",
									 -- x"59616248", x"2E222934", x"2F313F41", x"424C5158", x"6D52555C", x"57525938", x"39464B45", x"50505A57",
									 -- x"53431017", x"0F14110B", x"0D071006", x"7079656B", x"70573B48", x"5F666554", x"403F4039", x"3F322F3A",
									 -- x"39393443", x"3B3A3F37", x"3F453F43", x"463C4442", x"43383D44", x"484A4C4C", x"484D5654", x"4949463F",
									 -- x"424A4C4A", x"34473F45", x"43404140", x"494B656C", x"6A6B5446", x"56666760", x"6C635C57", x"655F5D54",
									 -- x"486E5D1C", x"46594559", x"3F5C6D4E", x"4139494D", x"4C484240", x"3B3E4C41", x"2C42454C", x"54574E50",
									 -- x"503F4E5D", x"3A33534F", x"6157554D", x"4E515064", x"3F495B6F", x"5035294E", x"6638343A", x"332D3435",
									 -- x"3D39464E", x"4E5D4A51", x"65705453", x"5C5A6760", x"5A65655F", x"61646469", x"5C60595D", x"5A5E7263",
									 -- x"5D9E9798", x"949B739A", x"B2A99778", x"9B9E9AAC", x"8A90859F", x"9874717B", x"91A1A9AA", x"9196927D",
									 -- x"8E6B5363", x"564B4E3F", x"68513642", x"3D7C3651", x"4B234C82", x"856B5251", x"64574F5C", x"62697279",
									 -- x"7B6A716D", x"74696E61", x"7266666C", x"63666A65", x"46536451", x"52555852", x"5C59616C", x"746F6683",
									 -- x"7E756A5A", x"8188837E", x"85897670", x"A4BA8F85", x"7F8F7C7B", x"897E8585", x"9A918285", x"88819792",
									 -- x"747D9399", x"95959AAB", x"A79B8484", x"8B8895AB", x"AD9D959C", x"889885A1", x"A6868A96", x"9B97878A",
									 -- x"7BA27F7F", x"799A7F87", x"7C99A092", x"8D808EA1", x"8B9C7A74", x"7C7C727F", x"776D7E92", x"596F6A5D",
									 -- x"62827E7B", x"7C5C685E", x"5D745249", x"5151675C", x"57425161", x"54595664", x"5A60725C", x"51566A66",
									 -- x"70597588", x"7C838578", x"7D699284", x"7E8A837C", x"7A95788D", x"6C6D7677", x"82694060", x"54645265",
									 -- x"60596B55", x"584F494E", x"54493845", x"41394B55", x"47565E5E", x"5E614654", x"7B7A616B", x"924B6686",
									 -- x"8585786A", x"CACBC4C0", x"C0BFBEC1", x"C5C2BCBD", x"BDBFC0C1", x"C4C7C7C6", x"C5C5C6C5", x"C5C5C6C7",
									 -- x"C4C3C1C2", x"C3C4C2C0", x"C2C2C0C0", x"C2C5C5C2", x"C0C1C2C3", x"C2C2C1C0", x"C4C5C4C0", x"BBB9B8B8",
									 -- x"B6BBC0C3", x"C4C4C6C8", x"C6C6C5C4", x"C2C2C4C6", x"CFD3D7D8", x"DADEE3E5", x"E8EAE8E5", x"E3E2DDD7",
									 -- x"D9D5D1D7", x"E6EEE6D8", x"D7DEE4DF", x"D2C5BEBD", x"B9A38267", x"5C5E5C57", x"554E455A", x"57665C48",
									 -- x"45394431", x"353C353B", x"3C3F3934", x"323A4036", x"2229223A", x"252E3334", x"323A3E3C", x"52484C4B",
									 -- x"514A515A", x"4E595356", x"53544B45", x"5446403C", x"3A393A3A", x"2F272527", x"2D333838", x"31313C38",
									 -- x"353C3D31", x"3838403D", x"3F3D4832", x"343C424B", x"48404640", x"47444447", x"494F4C3E", x"52544D52",
									 -- x"5E4F5185", x"5C58485C", x"4A235A60", x"5650484A", x"49494446", x"4F46383B", x"32143741", x"3A383D24",
									 -- x"344E3A47", x"504B4932", x"3E393849", x"463A2C35", x"454B5255", x"4E4C4E49", x"69626668", x"636B5A54",
									 -- x"78755D73", x"79706F4B", x"4966654B", x"626F566A", x"5E535758", x"55695D56", x"576B604D", x"555B527D",
									 -- x"56525D61", x"63586E5B", x"50565E68", x"5E555C59", x"5762615A", x"58585859", x"695F5851", x"5D676364",
									 -- x"769D8D7F", x"6E8994AB", x"C9A39B9C", x"BFAC9C51", x"898F649A", x"806D9374", x"9089869E", x"92A38879",
									 -- x"78665A74", x"4F70454B", x"4B6A2C1D", x"364A1F42", x"212A4130", x"47493E40", x"3D272A3A", x"4F5E595A",
									 -- x"5652525F", x"4F56575A", x"545A5856", x"484F555D", x"635D6E6D", x"68665E6F", x"5C60635D", x"5168478E",
									 -- x"6A466C65", x"719E6B78", x"7D76748A", x"8068667B", x"6A47635E", x"70785660", x"83776A6F", x"665A796B",
									 -- x"7D777677", x"6A6B746D", x"6E7E7872", x"716F7B8C", x"80787F7D", x"576F6E77", x"74685F72", x"736A756A",
									 -- x"5B5D8484", x"626A6B74", x"646C7369", x"5D5D7475", x"5B5C6E70", x"576A6676", x"7F6E635D", x"5C736C78",
									 -- x"B5785D69", x"50677250", x"484D4F6A", x"4E575854", x"4E4D524F", x"5F5C5756", x"575E6261", x"57545E62",
									 -- x"5C64686C", x"6C98716A", x"757C7C73", x"6A6F5C56", x"5D665062", x"5C886659", x"64716161", x"6F707173",
									 -- x"59545463", x"675B606D", x"64665D5E", x"58536265", x"625A5244", x"5259554F", x"3E5B5959", x"526E6269",
									 -- x"53506D54", x"6EB5B9CE", x"CEC7C9C2", x"BBBFC0BF", x"BDC1BDBD", x"C0C2C6C0", x"BFC2C5C3", x"C1C0C0BF",
									 -- x"C2C3C0BE", x"C1C1C0C3", x"C1C0BFC0", x"C2C3C1BF", x"C0C1C1C1", x"C0C1C2C3", x"C7C3C5C4", x"BCBBBDBA",
									 -- x"B9BDC2C4", x"C4C4C4C5", x"C6C6C8CA", x"CAC9C8C8", x"CBD4D9D6", x"D6DBDDDA", x"D6D3D9DF", x"DCD4CFCB",
									 -- x"CBCCD2D5", x"D9E3E2D3", x"D3C5C5D3", x"CCD3B787", x"887F6F45", x"4B644C48", x"3F343449", x"33393C3A",
									 -- x"3E363342", x"3D404B45", x"47434445", x"43474941", x"42463D3B", x"4C413E40", x"3F433D3B", x"464D4A47",
									 -- x"484B4551", x"4B484443", x"444C4442", x"40393F3F", x"332F393C", x"35312D32", x"37362E2C", x"2E2F332D",
									 -- x"30302F2E", x"2F323433", x"353B3741", x"3537413F", x"41414847", x"4E494C49", x"494E4B48", x"5F3F3B4E",
									 -- x"493D4243", x"48514538", x"36342E2F", x"3533181A", x"34213538", x"3C392A24", x"34352A2C", x"2A302F39",
									 -- x"41263153", x"38423D48", x"4346434E", x"524A504E", x"4B46465B", x"6A556E62", x"64646265", x"5B785444",
									 -- x"55595645", x"433B4044", x"45434333", x"4C363B45", x"4A564C42", x"38504949", x"4A504D47", x"3D453955",
									 -- x"34363B41", x"3A3E333F", x"484F5046", x"4B434543", x"44464C45", x"48474E4D", x"3A504549", x"444F522F",
									 -- x"8DB69977", x"5D8FA972", x"575592AB", x"9DAA9965", x"8A97838D", x"5A76754E", x"8FBA7C8D", x"B0708879",
									 -- x"72547B3A", x"4D683C38", x"37293228", x"4539678D", x"26413E39", x"3A363C3C", x"3C42443A", x"3C443E4B",
									 -- x"4D504744", x"4E4F4847", x"495B585E", x"655C677C", x"65626462", x"5D626660", x"5B6B5F64", x"5E6D6A7B",
									 -- x"6B727665", x"63636763", x"6A78695E", x"687B846C", x"6E736374", x"67845F57", x"5F68676F", x"69636458",
									 -- x"555B535D", x"85846A64", x"6571665E", x"5C555246", x"474F6449", x"65625E61", x"5A72695B", x"93656D75",
									 -- x"51415D5D", x"58715859", x"4145465A", x"635B5D54", x"61565969", x"656A6A72", x"62576F72", x"65648475",
									 -- x"585C4462", x"6B4B565F", x"78656669", x"6C5F5A78", x"66646550", x"415A5E57", x"4C5F6356", x"57595A67",
									 -- x"67616460", x"58635064", x"615A7368", x"6E6D8B82", x"797A75B0", x"8C7B7970", x"5D5B5C58", x"516B6C65",
									 -- x"6063646B", x"6E6C6F6A", x"5B6D736E", x"74766C6A", x"73818778", x"84846E58", x"5E675F5B", x"474E4B61",
									 -- x"6D6B6E6D", x"67677386", x"9E9DA3B5", x"C3C5C5C7", x"CBC9C1C3", x"C4C1C1BC", x"C4C0BDBD", x"C1C3C3C2",
									 -- x"C0C2C1BF", x"C0BEBDC0", x"C1C2C3C3", x"C1BEBCBA", x"BEBDBDBF", x"C1C2C3C3", x"C6C7C2C2", x"BDBDB9BB",
									 -- x"C4C5C6C6", x"C6C6C5C5", x"C7C6C5C4", x"C4C5C6C7", x"C4CACFD1", x"D1D2D4D5", x"CCCCCCC9", x"C4C6C7C4",
									 -- x"C1C0C3C5", x"C6CCC9BC", x"CDD4C3B2", x"9A784938", x"6365674E", x"433F2E3C", x"40433B3C", x"3C403F42",
									 -- x"3F485B54", x"42524F4D", x"56515253", x"4B43454B", x"424A443A", x"413D4850", x"4E555859", x"5C5E5B58",
									 -- x"44413F3C", x"40373D39", x"42403B40", x"42343534", x"31333937", x"302F3133", x"2B313232", x"3739403B",
									 -- x"3B393839", x"3B3C3A39", x"41423E42", x"3E414747", x"4B48444A", x"4D524B46", x"43443D41", x"2F212E29",
									 -- x"27233034", x"29212436", x"191F3331", x"1E323C37", x"3A463D2C", x"3B4B584E", x"54535F67", x"51575F5C",
									 -- x"535B4E64", x"59757A8C", x"6967585F", x"575B4C73", x"5C69666B", x"544E524D", x"5833353B", x"4D4F464B",
									 -- x"483D3F47", x"40373639", x"39393745", x"46433B43", x"40494145", x"3F54484B", x"4747414E", x"454A4B42",
									 -- x"4A494C4C", x"41433F4C", x"3B324B48", x"494B474D", x"52475058", x"48485252", x"5252554B", x"4C574E33",
									 -- x"92876668", x"82B69894", x"7D2B2F76", x"B39D9D96", x"88837A89", x"877F7454", x"728C9D93", x"6F769840",
									 -- x"58987F40", x"30313329", x"34363A36", x"423C3E41", x"45372E34", x"42382B3A", x"383A3539", x"383F3C35",
									 -- x"46484244", x"3F4C4D4D", x"4E554E60", x"6057546F", x"72686560", x"56555A59", x"5966595D", x"63604E5B",
									 -- x"594D655E", x"515A5D5F", x"5F5C685D", x"535D554A", x"689D684A", x"404E555F", x"57595A6C", x"5C7A655A",
									 -- x"4B565541", x"5D5A6967", x"5770675C", x"68725F5C", x"63636461", x"686B6660", x"6170797F", x"9B6A6377",
									 -- x"60705965", x"70786A66", x"70607D7A", x"5B63775F", x"615D4362", x"73575867", x"6C79888F", x"937B7878",
									 -- x"6B685D7D", x"897F8668", x"82706F60", x"5D627564", x"64685E5A", x"6B647086", x"775E6664", x"6966596A",
									 -- x"805E6B5C", x"64616864", x"5B58606D", x"7959698A", x"905C7666", x"616E756D", x"6B6D7975", x"6B685E6D",
									 -- x"78767272", x"70767D72", x"717A7E78", x"84806872", x"787C827C", x"82787A8D", x"857A7989", x"8E8B726B",
									 -- x"73706272", x"786B6F67", x"6C6D6563", x"6E7C8A92", x"98999CAE", x"BDC2C8C8", x"CBC6C4C6", x"C7C3C0BF",
									 -- x"BFC3C3C1", x"C1BFBDC0", x"BEBFBFBB", x"B7B6B9BC", x"BAB9B9BB", x"BDBFBEBD", x"BCC3BCBE", x"BEC1BAC0",
									 -- x"BDBCBBBC", x"BEBFBFBF", x"C4C3C1BF", x"BEBEBFBF", x"C3C4C7CA", x"C8C4C3C5", x"C7C3C4C6", x"C6C7C6C1",
									 -- x"CDC8C6C4", x"BFBCB7AD", x"95866955", x"47434654", x"41454A4A", x"4D4A4758", x"444C4E46", x"453F4146",
									 -- x"4B518959", x"4B50494F", x"4E4E4F4F", x"4C454751", x"494C4E4E", x"544D5555", x"5351514F", x"4A474642",
									 -- x"3C3A3631", x"39384442", x"40352F2F", x"39323938", x"343B3C3A", x"38393A34", x"3A3A3C3D", x"3F333B3C",
									 -- x"37383B3E", x"3E3C3D40", x"38383C3B", x"403A2F2B", x"41404A41", x"4A404947", x"44483847", x"443F5049",
									 -- x"5053544A", x"494F4F54", x"49584944", x"565D5169", x"6E805947", x"7A795F5E", x"5A555F61", x"494B4E40",
									 -- x"38484D56", x"594B5255", x"4F3D4B56", x"4E52463A", x"4249464D", x"3E4A3F39", x"43434842", x"48354E4A",
									 -- x"42363D54", x"4845423F", x"403F3F40", x"3F454641", x"3E464141", x"2F383345", x"473E433B", x"3D4B3F47",
									 -- x"453E4044", x"41413938", x"3E384D41", x"3B4C504B", x"4250494D", x"4B44384A", x"47495646", x"3E3F4541",
									 -- x"60384466", x"78957E97", x"ACADA18D", x"9292A87C", x"7CA1715C", x"82427A5E", x"4A79888C", x"7E737D5D",
									 -- x"4E704A44", x"4A3D3E45", x"3B3B393C", x"42403B3D", x"3C334C45", x"40564D3F", x"41344834", x"4E4F4644",
									 -- x"43413E4C", x"475A5141", x"57504A55", x"5C56526D", x"645A534E", x"4E58584B", x"6653535B", x"5F6D705B",
									 -- x"5A64645F", x"5A5A5A63", x"5C4C4D63", x"504E6D53", x"4D35564C", x"5C605F60", x"47566860", x"60565855",
									 -- x"61536266", x"4F636355", x"62725E41", x"5961506A", x"685C5A61", x"4C535F53", x"63637066", x"5861674D",
									 -- x"696D6062", x"6262644E", x"4B4B565E", x"554F6663", x"6668645B", x"59525457", x"525B6671", x"6C575F70",
									 -- x"6B747F7B", x"76757679", x"87706D6C", x"4B6D6664", x"42656763", x"5D6B6359", x"57496564", x"5E676956",
									 -- x"65653D6E", x"727A655C", x"727C6467", x"5E6B696D", x"586B7463", x"7F93826F", x"8591796D", x"674F555A",
									 -- x"6E63636E", x"71788786", x"85847E7A", x"837E717D", x"75736C5E", x"6C6E6E78", x"77767A75", x"6E72757A",
									 -- x"74777B79", x"76726B66", x"7670736B", x"666D6967", x"65625D66", x"717A878B", x"989BA4AD", x"B0B0B6C0",
									 -- x"BFC3C4C6", x"CACACACD", x"CCCCCAC5", x"C0BFC1C5", x"BCBCBCBD", x"BEBEBDBD", x"BFC4BFC2", x"BCC0BBBD",
									 -- x"BCBBBBBB", x"BCBDBEBF", x"BBBDBFBF", x"C1C2C2C1", x"C2C3C6CC", x"CECDCCCC", x"C4B2AEB7", x"B6ABA29E",
									 -- x"988F8780", x"756A625D", x"5E54555F", x"5F656B6A", x"68655855", x"5C5D5955", x"5F4E565C", x"58545653",
									 -- x"5B5F4A51", x"4C566255", x"6065615B", x"60615D5D", x"645A5A5E", x"5A494A45", x"39313339", x"3B404440",
									 -- x"3F42373B", x"39444949", x"4D494940", x"484A5147", x"42453D3C", x"40413E34", x"3C3B3C35", x"372D3939",
									 -- x"3D404544", x"3C363A42", x"4641463D", x"4A494143", x"4C4F5C4D", x"4F3F4C4F", x"5C503F4A", x"6253564F",
									 -- x"697A7457", x"4E555552", x"48414D5E", x"50505251", x"473B4C4F", x"5C594544", x"423F3C40", x"474C402F",
									 -- x"32334A50", x"4D394A46", x"4A4B413D", x"403B453C", x"443E4044", x"47413F3E", x"433F3E42", x"433D4B4E",
									 -- x"47474C52", x"474A463C", x"42413F33", x"393B423F", x"3F3A3432", x"31363139", x"38264138", x"323D2C33",
									 -- x"2315141A", x"29374243", x"383D3A34", x"2F3A4B3C", x"26383F3F", x"3B423E37", x"3F372F37", x"3A2D280C",
									 -- x"77412C2F", x"43413F4D", x"486995A4", x"5B588670", x"44534927", x"37494351", x"3E2F617E", x"614F3F4A",
									 -- x"483E4040", x"464B4745", x"42464F4A", x"4C434749", x"4C434B42", x"48584F53", x"496B585A", x"4D424756",
									 -- x"55575554", x"4D5A5E5B", x"6154584A", x"5A50505D", x"59514F4E", x"515B5B4C", x"41535C4A", x"5455574F",
									 -- x"66595E57", x"56543763", x"54414850", x"464D5B5B", x"52515258", x"4F61525F", x"67595D5B", x"5A4E4749",
									 -- x"494D735D", x"58695E5B", x"54638872", x"5C5F7266", x"5F666564", x"6C665F5F", x"626C6665", x"69716E64",
									 -- x"5462685F", x"6B5D7863", x"62736A45", x"58684452", x"5E5A6659", x"56555658", x"5E64645D", x"4D4B5758",
									 -- x"504C6366", x"50444C46", x"696A6872", x"6A5E6964", x"4640695F", x"5C666F44", x"65616169", x"624A5B5A",
									 -- x"687C536D", x"707A6B65", x"796F6170", x"727A7181", x"8A7779B0", x"6F516F62", x"5A65716A", x"6F60565E",
									 -- x"6A626675", x"726F7876", x"7C858180", x"8387897F", x"7C78756A", x"716A6164", x"635F635D", x"6167635C",
									 -- x"7267695D", x"5864799B", x"8A5D6364", x"606A6369", x"636A6B6E", x"6E68655B", x"6767696A", x"66646E7B",
									 -- x"7477787C", x"8487888A", x"979DA5AC", x"B1B5B7B8", x"BBBEC0C0", x"BFBEBFC1", x"C1C0C2C6", x"BDC4C5C1",
									 -- x"C4C4C3C1", x"BDBABABA", x"B5B5B3AC", x"A6A09A95", x"99999795", x"95938E87", x"87746C71", x"6E646162",
									 -- x"635F5D60", x"63616267", x"686B6C6B", x"6C696868", x"60666061", x"6565655E", x"625E6965", x"4D495265",
									 -- x"63646C6D", x"7670756C", x"7A7D746C", x"6E6C625C", x"5C524E47", x"3C323F3E", x"3E393F47", x"4A4D504C",
									 -- x"494E464C", x"4C555755", x"56525345", x"4348504B", x"43443B3A", x"42454544", x"3D454235", x"3639433B",
									 -- x"41424545", x"413E434B", x"504A4D41", x"4B4C484E", x"42463E4A", x"414D4447", x"513A3C46", x"5455544D",
									 -- x"4B545045", x"3C323138", x"343E3532", x"31363948", x"41364F46", x"3B3C3B3C", x"3B39373A", x"48493823",
									 -- x"20232F37", x"2432353D", x"3F42344B", x"40403B3B", x"3C40443E", x"35162833", x"3E313B38", x"37483B42",
									 -- x"4046453B", x"4147473E", x"3540373A", x"3D3C333D", x"2B2C322A", x"32302F31", x"292D2B30", x"382D252B",
									 -- x"2F2A2D29", x"2F2B3331", x"2C302735", x"3A343D3D", x"39484E42", x"464D4D3F", x"46453B3C", x"28222E31",
									 -- x"412B3939", x"261B3129", x"314A343A", x"35443C44", x"463A4138", x"3B394037", x"4D4A3E4A", x"38344042",
									 -- x"3D3D423E", x"303B483A", x"2C3B453A", x"3B42463B", x"453D4A45", x"2D3A5049", x"4A50434B", x"444B4747",
									 -- x"4E514F44", x"4A443F3A", x"3E38463E", x"524D4E56", x"544E4F4E", x"45444948", x"4A656C50", x"5F524E4C",
									 -- x"55534E51", x"46484848", x"35494D4A", x"504C4C61", x"3D485C62", x"5F705C5A", x"72515E6E", x"665D5766",
									 -- x"4D354D50", x"3C3E4E56", x"5B576168", x"5749595C", x"645B5D53", x"51605D5D", x"55625C61", x"615F6B5D",
									 -- x"63665B58", x"4E428E6A", x"5F755956", x"6775666A", x"6F89807A", x"7C616769", x"5B6E6B68", x"727F7A65",
									 -- x"5B6B5E70", x"89707471", x"69698284", x"9999826D", x"6E6D6A69", x"62849171", x"687A6768", x"7F6A6873",
									 -- x"686E7464", x"5463675F", x"5C696D55", x"80876B66", x"7066596D", x"63667361", x"766E5C72", x"81677067",
									 -- x"54585E65", x"63646B65", x"666C6668", x"635B5E50", x"5E555D5B", x"55434456", x"51525958", x"58595960",
									 -- x"5F5B595E", x"5F5F6B77", x"6C4A585C", x"58615756", x"5A5F5B59", x"5B5F6764", x"64616061", x"6061656B",
									 -- x"60636364", x"6969686B", x"5F616468", x"6A6A6968", x"6366696A", x"68696C6F", x"76737575", x"757B7F79",
									 -- x"797B7B78", x"726E6C6D", x"68696763", x"6061605D", x"60636464", x"676A6964", x"66646563", x"5D5E6364",
									 -- x"64646264", x"68666870", x"66636C6B", x"676A6F61", x"5D60646A", x"68626567", x"67675F5B", x"6A74646E",
									 -- x"6A755969", x"6069665B", x"5A585453", x"51494446", x"4B4C4D46", x"464A574C", x"46474A49", x"44444748",
									 -- x"4A4A4B49", x"524C5148", x"4D484F4E", x"44494D50", x"46494A43", x"47484148", x"4B4A4549", x"46404244",
									 -- x"4F4D4B4D", x"50535555", x"4341423A", x"3B383437", x"3A3A303F", x"3D4C4444", x"44454342", x"3C4A3C46",
									 -- x"3D39343F", x"4337302E", x"4144373D", x"42433A38", x"3C40322E", x"423C3A3C", x"3C353C3B", x"36343424",
									 -- x"161A2633", x"33392E41", x"412E363F", x"36473A2D", x"2A363130", x"2719252E", x"3441453C", x"32303932",
									 -- x"38383329", x"3B3F423F", x"30464133", x"3C3A2D2B", x"252F3D2D", x"2C262C34", x"3233373C", x"3533363F",
									 -- x"40382E20", x"30293737", x"35353336", x"3A3D333C", x"444D4637", x"47413D41", x"42374248", x"3F4A3D41",
									 -- x"3A443F3B", x"42463748", x"3F4A4647", x"45473D45", x"404A3D46", x"3C3D3B51", x"4842443D", x"3247453C",
									 -- x"3E403445", x"404A4647", x"4B4C4442", x"3B474238", x"3B454651", x"42273F61", x"52316748", x"3E47464B",
									 -- x"463B3027", x"464A4F4F", x"49434148", x"47464250", x"4C4C4B40", x"3D4B5144", x"413D443C", x"50434238",
									 -- x"4C4C5446", x"4351413F", x"4754505A", x"514A625B", x"5F50557E", x"3844493E", x"4B6A3C30", x"47526140",
									 -- x"3D412B56", x"5344506B", x"5F474370", x"605D635F", x"5B464855", x"59795C45", x"7B565475", x"604B6C5F",
									 -- x"6171564D", x"4D4B5C5B", x"625B5F6B", x"67614A68", x"66696669", x"6B606562", x"6B61646E", x"6F6F786C",
									 -- x"65585D59", x"68655C52", x"53645A59", x"515F776C", x"8B90796F", x"7F52676E", x"6B5A616C", x"6D604D5A",
									 -- x"5C5C4B67", x"5B5C5647", x"5C5E5F56", x"5D65515B", x"585F5153", x"57565252", x"805E4A43", x"525D5C63",
									 -- x"5F65615C", x"585A5F5A", x"5A5A5861", x"6B6A6C73", x"605C665F", x"60605D53", x"50555959", x"59564F59",
									 -- x"545F6061", x"5C575B58", x"6161645E", x"5C605B52", x"57595556", x"58585D5A", x"5A585759", x"5C5D5C5A",
									 -- x"5D626361", x"615D5B5E", x"61605F5E", x"5F616364", x"65676969", x"68696B6D", x"6C6A6255", x"68676664",
									 -- x"686A6B6A", x"69676565", x"6A6C6965", x"64676867", x"64656868", x"66646567", x"5F646968", x"6161625E",
									 -- x"666A6869", x"6C69686F", x"74677477", x"75787D65", x"6F65666A", x"6A676669", x"69666355", x"67644F53",
									 -- x"50576656", x"52504E54", x"524F5052", x"4F4D4F51", x"46494E50", x"56555B50", x"545A5A56", x"565A5F64",
									 -- x"6F6B6966", x"695D5D54", x"47495964", x"575F5652", x"4D505443", x"474C393F", x"44413C51", x"49403D48",
									 -- x"4A4A4642", x"41423D37", x"41403939", x"34384143", x"3E3B3B35", x"38363A3A", x"35413A3A", x"343F333E",
									 -- x"3A414041", x"39313229", x"3D3F3539", x"33383F3D", x"4333343C", x"3D373D30", x"312F3736", x"393A4647",
									 -- x"3A2B2E32", x"37282A33", x"2E3B3E27", x"33332427", x"2C322C2E", x"2F322C31", x"3B352936", x"382C3E3C",
									 -- x"3C3A3831", x"30333633", x"39423E2B", x"35342E24", x"37363532", x"373C3638", x"33234854", x"27394736",
									 -- x"3F3C342B", x"4A3E443D", x"3A3E3930", x"28363331", x"2F222C35", x"2E2E3730", x"432F3735", x"38463732",
									 -- x"413E3E3F", x"3A493D40", x"463E4148", x"4B3F3C43", x"404B4338", x"4D453A48", x"42453B43", x"3E3C453E",
									 -- x"4349393F", x"454E4146", x"443F434F", x"4A4A4744", x"424B3E37", x"2E2F4544", x"3C34404A", x"3B464E48",
									 -- x"3E3E4440", x"453E464C", x"4644363D", x"363B3F48", x"4C484444", x"51676449", x"3D4E5750", x"6549414F",
									 -- x"56534656", x"5D41434F", x"65445355", x"3C41473C", x"6B4B543F", x"4C4F3B38", x"546F293E", x"3A2A4F56",
									 -- x"475B5E63", x"594C6A5C", x"475C5852", x"47504E50", x"40555250", x"525D556F", x"565A4D58", x"5E5B5F5A",
									 -- x"524E6770", x"667C5F58", x"51646B78", x"77686E6F", x"814A4E6A", x"6661595C", x"614E5C60", x"4F4A6B6B",
									 -- x"5549564A", x"64644D4A", x"595E5D47", x"5B5E6259", x"6A76716E", x"71667076", x"816F7A70", x"576D635A",
									 -- x"6157414A", x"5A4C4E37", x"52575867", x"404F647C", x"655F424F", x"4E4E4F5C", x"5864574F", x"52524D4E",
									 -- x"4C514A48", x"49494E4E", x"545A5549", x"5861555E", x"584C5B60", x"5F5B6061", x"6168625E", x"62695F66",
									 -- x"5E5D6768", x"6A6A6161", x"5B645154", x"60595954", x"625D565A", x"5B575A5A", x"5C5B5958", x"5A5E605F",
									 -- x"5A636766", x"635F5E64", x"63646565", x"65656566", x"6A6A6968", x"67676768", x"60635444", x"6D6B676D",
									 -- x"63646566", x"68686766", x"6B6D6D6A", x"6B6F716F", x"66676B6E", x"6962656E", x"736F737A", x"79757372",
									 -- x"73797774", x"766F6B71", x"70726C62", x"726C686A", x"665C5D5C", x"5C605D5B", x"5C46544C", x"59535154",
									 -- x"575E5758", x"5A4E5857", x"5A585751", x"4D53554A", x"5250555B", x"5E556773", x"6B726D65", x"65625A56",
									 -- x"53534B56", x"52524D4C", x"46454543", x"314B453F", x"3C3A3E2C", x"3F5A4B53", x"3F4E484E", x"4047403C",
									 -- x"3E454741", x"3D3C3934", x"363A3540", x"36373C36", x"3B3C3638", x"31383A40", x"422F3546", x"3C3D4835",
									 -- x"3B414140", x"332E3832", x"344F4031", x"2F40453A", x"432F372F", x"363D332D", x"2B332D26", x"3C332D38",
									 -- x"3C2B242F", x"212D3F2F", x"31341F2C", x"29343533", x"3439453D", x"39352D41", x"352A403A", x"41634544",
									 -- x"3B434A46", x"303B443E", x"483A2B46", x"3B3E3240", x"3B3A353D", x"383E2B2C", x"1E3D262E", x"2B2E322D",
									 -- x"34383024", x"45374040", x"33382C37", x"272B3F34", x"33383E4C", x"47433A3A", x"4740423E", x"3F3D4236",
									 -- x"383B4244", x"3C3E483C", x"403E4B54", x"403D4F4B", x"4F444551", x"464F4845", x"303B4645", x"43423B3B",
									 -- x"42371B2E", x"43334745", x"3B3F5146", x"423A4843", x"48574A45", x"4A434753", x"414D4242", x"443E4047",
									 -- x"3B39454B", x"413D474D", x"4F54463E", x"3B3E473E", x"452F314B", x"5955493D", x"41405148", x"44374544",
									 -- x"3F3B3E40", x"3C394B3D", x"38373951", x"4F3A3E3F", x"3A5B5343", x"814E4449", x"5234545F", x"675D7F60",
									 -- x"67574B56", x"4B525261", x"55455748", x"433D494A", x"61464D4A", x"31314F41", x"474F474F", x"50514E63",
									 -- x"5D4C5D64", x"576A6152", x"594F6268", x"6353665A", x"5557556E", x"62556067", x"5C7A8971", x"7374857A",
									 -- x"6262595F", x"5C446959", x"5494806B", x"686C6A80", x"C7788F87", x"7D87938D", x"99917D83", x"7A76606B",
									 -- x"645E8D54", x"43656650", x"666C6162", x"665E756D", x"625C6563", x"615C5669", x"67655656", x"6E775863",
									 -- x"4A52504E", x"53504D55", x"6062565A", x"6151474E", x"4C524947", x"4446424A", x"3C484F4F", x"53595955",
									 -- x"625F5D62", x"665F595D", x"5B5A4445", x"50534955", x"55545754", x"48534F54", x"634E4C57", x"57575F63",
									 -- x"59626866", x"63656767", x"6A6B6767", x"6265657B", x"6D6A6066", x"57646262", x"564F4C46", x"57585559",
									 -- x"5D575D5C", x"5A615E59", x"605E5F5E", x"5D5F605B", x"5C5A5762", x"5E615F67", x"68657066", x"63685F65",
									 -- x"65646568", x"68656363", x"5B5D5A5D", x"5F5F615D", x"5E595654", x"53575954", x"52585058", x"5A5A6456",
									 -- x"584D5C62", x"5C565E50", x"4F4F5455", x"50545955", x"594D5354", x"414B5053", x"4C565051", x"50524748",
									 -- x"4149484D", x"4D524C4D", x"4844474B", x"4442463D", x"372B4442", x"41353B3E", x"332B353A", x"362F2D34",
									 -- x"33313833", x"38333A3A", x"372F3C3C", x"3C3F373B", x"37323636", x"33373233", x"2A293838", x"39323331",
									 -- x"3C3C3632", x"3B373426", x"2A313130", x"223F3D39", x"3B3D2B35", x"3C323730", x"2732232D", x"322E2932",
									 -- x"38382F2C", x"3236383B", x"39403C3C", x"3B433E3C", x"403F453E", x"3E3B4342", x"46404540", x"433A3739",
									 -- x"38343724", x"3E493B42", x"4546463B", x"443F483C", x"373C322F", x"3F49323A", x"354A422D", x"43394042",
									 -- x"3A3C5736", x"302F484F", x"42393E48", x"3D465C4E", x"595D4351", x"483F3A3C", x"42415044", x"3C4A4644",
									 -- x"49424D4B", x"46504A4F", x"4D475D58", x"495D4C49", x"4E474649", x"4C51514B", x"4A414046", x"4A474748",
									 -- x"4545493E", x"515D5244", x"4B485D55", x"39556364", x"4D505256", x"4F5F5152", x"614C454A", x"4F444D4A",
									 -- x"4F574E53", x"5747454F", x"4B674F40", x"47493C3E", x"43461744", x"45454341", x"403B4220", x"3B3E3B3F",
									 -- x"2E3C3D37", x"44434736", x"3C4A475C", x"4A425447", x"5153515D", x"5E4C604E", x"5281916B", x"5B594249",
									 -- x"5B4E2D45", x"4C78394D", x"394A4E55", x"4E414B44", x"4F3A4447", x"4C50372B", x"424B3A4F", x"59485154",
									 -- x"5447544F", x"3F506356", x"50515F60", x"57525D48", x"63875869", x"5C585975", x"65786F50", x"677C4F63",
									 -- x"575C6353", x"5E62716E", x"697C676C", x"6A606666", x"97706150", x"6D8C8B87", x"74707475", x"6B5B6966",
									 -- x"5E607791", x"766A6E69", x"66636262", x"5A5E595E", x"57606365", x"68636269", x"67676B4D", x"696C5E76",
									 -- x"4E575B5A", x"57504F58", x"54564C51", x"50474A5B", x"4C3F373E", x"3C494B45", x"444E5356", x"5A595454",
									 -- x"53554F4D", x"524F4C51", x"4C41342F", x"35323135", x"3629354A", x"44413331", x"403B3A4A", x"5D615E61",
									 -- x"5E626462", x"61636463", x"6562605B", x"55555460", x"57534E51", x"51585248", x"52545752", x"59575155",
									 -- x"565E5E58", x"5C595363", x"5C5D5F5C", x"57595E5D", x"5D5F5E66", x"63645C5B", x"63666B5C", x"57605956",
									 -- x"575B5C58", x"55555757", x"535B5C5E", x"5A555A5A", x"5F575251", x"51565B5B", x"685C5E5B", x"5A5C5455",
									 -- x"4C525252", x"5156564D", x"504F4F4D", x"4C50504A", x"424E3539", x"45404244", x"49484741", x"4F47413A",
									 -- x"3637425A", x"4D474B49", x"4F49454D", x"45464848", x"4842443B", x"3E494839", x"40373133", x"32433E3C",
									 -- x"3C373645", x"48453A3B", x"3E443F35", x"3C40333E", x"2F2E3639", x"392F2D32", x"322D2A2F", x"262C3039",
									 -- x"2C394031", x"38342330", x"2A293329", x"3D3C453F", x"2F2F2531", x"33272D27", x"33272833", x"3633352C",
									 -- x"40353849", x"513F4239", x"3C303039", x"303F473E", x"3640422E", x"313B4743", x"46444044", x"4945444A",
									 -- x"4947434C", x"54563842", x"4A504B31", x"3F4C6255", x"41393942", x"4E5A4E40", x"536C4E4A", x"3D304D44",
									 -- x"3B584B45", x"474B473F", x"5050443F", x"3D3D423C", x"363E3E50", x"47376046", x"59454052", x"4653414C",
									 -- x"4C474C3E", x"484E474A", x"534B4E46", x"414F4249", x"484A4A47", x"4F5F6050", x"52615656", x"54574B49",
									 -- x"535A5B51", x"474D474F", x"4B434E50", x"465B3C4C", x"42425041", x"494C4A39", x"4B3B3A50", x"3B434D4A",
									 -- x"4F505B40", x"43454C4E", x"53435658", x"555C5454", x"44484858", x"604C5155", x"4F3C4838", x"533E4C58",
									 -- x"504A4E48", x"59765A4B", x"443E485A", x"4A586155", x"555C5256", x"5C3E363D", x"2B445D5E", x"5D3E474B",
									 -- x"42415652", x"5C55514D", x"5F5B4B3E", x"54574F50", x"53545256", x"56524F41", x"5345444E", x"5A57683C",
									 -- x"49504E56", x"4F55515C", x"424F6159", x"5E525C69", x"56834F4B", x"514F5864", x"7169635A", x"5A49514F",
									 -- x"4B495C6F", x"5D60756C", x"736A6B65", x"595D6069", x"5F6A7C7E", x"6D7B7A72", x"7365515B", x"565A6163",
									 -- x"616A769F", x"A66B6C5D", x"5A606361", x"56566162", x"69685D54", x"566A6471", x"706C6D86", x"61536355",
									 -- x"54565A58", x"4C454D58", x"52524A52", x"44393844", x"303F403C", x"3A525549", x"4454554F", x"504F4D55",
									 -- x"4B4E443E", x"494E4B4F", x"40363631", x"332A2C26", x"222C353E", x"37251E3D", x"312B313A", x"404D5755",
									 -- x"5C5D5D5E", x"5F616160", x"625E6560", x"5F5F5E5E", x"5D5E615F", x"63605E57", x"5E65665F", x"5C62646F",
									 -- x"5D615E5B", x"635F5969", x"64646562", x"5C5E6363", x"67696566", x"6467605A", x"51575850", x"50595A55",
									 -- x"515A5F5A", x"595F6667", x"60646264", x"625E615F", x"615A595C", x"5B5B5D5D", x"615E6154", x"525C534F",
									 -- x"50654C50", x"5C574846", x"4446413B", x"3F433F39", x"403A4C43", x"3E484850", x"45484248", x"45494045",
									 -- x"434B434A", x"4B484543", x"4341413F", x"40414240", x"3C3D4146", x"473F4546", x"42383448", x"46514141",
									 -- x"3841343E", x"39382734", x"4B382C42", x"3D434129", x"2F323534", x"3C2C3034", x"36322D31", x"3332352D",
									 -- x"34262F2D", x"23313832", x"252C2D38", x"2E3C3B2F", x"25302A30", x"3020232D", x"28353232", x"34392F3B",
									 -- x"3C313641", x"493F4E37", x"3A38352F", x"22373E2E", x"3D3D352D", x"3E484D4D", x"524E4042", x"51474F56",
									 -- x"565C515B", x"4F4E4866", x"604F4A5C", x"604D4E57", x"51575459", x"6B624E3C", x"4769393D", x"5A4C4538",
									 -- x"363B2742", x"4855473D", x"4A474337", x"232C4442", x"3940493D", x"3E37514B", x"5A494845", x"43494142",
									 -- x"3F454C48", x"4F4E414B", x"454B4B4B", x"4F534C5A", x"4B464547", x"4D545147", x"42534D50", x"5A4A4854",
									 -- x"59536154", x"5133394A", x"50554F54", x"60505555", x"65564F50", x"4558616B", x"5D564B5E", x"59605D5D",
									 -- x"54586764", x"5E576B59", x"635D576D", x"87829390", x"998C8379", x"696C94A8", x"8579785B", x"5E65535E",
									 -- x"6B656766", x"5F56525A", x"7481676B", x"7F857185", x"6B6C6F6D", x"7F867962", x"78626F63", x"566D6D6D",
									 -- x"66605F80", x"6D5E5E4C", x"655D6574", x"5C5E5A5A", x"58625F5E", x"5B5E6059", x"614B434B", x"5A536956",
									 -- x"5360584A", x"47565247", x"55575A53", x"5953546E", x"56525157", x"5649624F", x"5957606D", x"6E4B5B57",
									 -- x"59566472", x"77566475", x"6D5B605B", x"5C615E69", x"86736F81", x"6F6C736D", x"5E524450", x"6F5B5159",
									 -- x"6B776752", x"4E685E5D", x"33464C3E", x"4C5B505D", x"5C555856", x"52564961", x"6574677C", x"6B555058",
									 -- x"544E5354", x"4744515A", x"4E48424F", x"3E312826", x"2E50504F", x"626E5446", x"47585347", x"4D4F4A4D",
									 -- x"43423532", x"43494446", x"413F4240", x"433C3B3B", x"3D3B3F3C", x"2D2A3139", x"112D3231", x"3E3E3944",
									 -- x"4F4F5152", x"53535353", x"5A545F58", x"5A5C605A", x"5E5D5E5B", x"59535355", x"545A5851", x"454D4C55",
									 -- x"57515756", x"52575959", x"64616160", x"5D5F605D", x"5C5C5A5A", x"5B5D5A57", x"57575357", x"57555959",
									 -- x"575D605D", x"5C5F6262", x"64635D5E", x"5F5C605F", x"625B5B5F", x"5D585656", x"52595759", x"51464E56",
									 -- x"5835434C", x"44473B4F", x"444C4841", x"464A4643", x"42423B3A", x"48414849", x"4F4A3744", x"3C483B3F",
									 -- x"4546423D", x"3E454343", x"373A4131", x"3D3A3629", x"2F404841", x"463A4135", x"2B242739", x"3030252E",
									 -- x"24202C33", x"1E2F3C2F", x"3934413B", x"2B371C2E", x"342F2E31", x"432D333D", x"33332F37", x"2F3E393A",
									 -- x"363D2E37", x"39363F37", x"3239353A", x"31333634", x"39312E34", x"3330312C", x"2C343B31", x"30414144",
									 -- x"3D3A3C3C", x"3F445143", x"394A453D", x"3D484546", x"49443A3C", x"4E4E494C", x"524E413F", x"58393B35",
									 -- x"28494640", x"3F484132", x"45483538", x"364A4942", x"45504034", x"3E2E2A27", x"3D312A31", x"524B4959",
									 -- x"433A2D36", x"53543644", x"4A414546", x"3E4C5641", x"3D474439", x"3F494656", x"4E515E51", x"595F5D52",
									 -- x"524E4E54", x"50524D5F", x"444F4F53", x"59554F50", x"554D4A4A", x"443F3A35", x"43474154", x"614E4F5C",
									 -- x"565E684B", x"5A596358", x"57575D5E", x"68637972", x"6B625B76", x"55625C69", x"57637261", x"59677E66",
									 -- x"624E6E8E", x"6E5A5963", x"6273A29E", x"7661625B", x"5A4E5137", x"3D4D2639", x"3F322B38", x"383B3839",
									 -- x"374C4238", x"56647642", x"53554867", x"5E606E73", x"635E6B4F", x"8F8C8954", x"646D6668", x"675A5968",
									 -- x"576C5288", x"6E6E766F", x"665D5C76", x"74695B55", x"5B555148", x"4053444A", x"60584F5F", x"604C4A52",
									 -- x"5D644A3E", x"4948495E", x"4F494955", x"4B4E4347", x"58484857", x"45494F60", x"56484846", x"474D4D4F",
									 -- x"50596B58", x"58585D4A", x"4856544F", x"584E4B5C", x"61687572", x"6E6B715C", x"52535252", x"5F4B464F",
									 -- x"46504535", x"4C4B4A49", x"3F3B4760", x"474B635F", x"47475355", x"5A535369", x"5E646B6D", x"6C606862",
									 -- x"42383F48", x"41414949", x"453E3D4B", x"423D3B36", x"43524947", x"4A453F56", x"464E4848", x"56544543",
									 -- x"403D3435", x"41423D41", x"464E4544", x"48494653", x"545F5044", x"514D4143", x"4C525752", x"4B4E4F45",
									 -- x"4D4E4F4D", x"4B4B4E51", x"57515A52", x"54585E59", x"645B5354", x"4C474343", x"40474F54", x"4F574F50",
									 -- x"50556057", x"4C525656", x"5655595A", x"55545553", x"51515659", x"5C585756", x"5A59565B", x"5B56595A",
									 -- x"58565658", x"5A595552", x"565A5758", x"524E565C", x"534A484A", x"47434445", x"4C4D4341", x"45434344",
									 -- x"3E363638", x"43454131", x"38454640", x"41444345", x"4B464D52", x"4C405152", x"45383129", x"28232729",
									 -- x"26163F4D", x"3D444B4A", x"49494C42", x"46483C34", x"504E3E3B", x"3F342915", x"2D323E3D", x"33333133",
									 -- x"373C3B34", x"48453D33", x"3C4F3B3F", x"34383C3A", x"2D383A2B", x"3B363D3C", x"40273834", x"3A3E323D",
									 -- x"2A39343A", x"3E364043", x"40423735", x"39343643", x"4A37464C", x"39404C40", x"40444B33", x"413A3B48",
									 -- x"4344464B", x"45453F49", x"3D403D4C", x"534D475A", x"37454848", x"4A41312E", x"3C3A2933", x"4F404341",
									 -- x"4D4B3A47", x"463B3D46", x"3435374A", x"4C464446", x"3E3D3B33", x"2B273C36", x"3A3F4835", x"444D3F49",
									 -- x"4B384745", x"43474134", x"3A494E46", x"44443E3B", x"3246364D", x"4D4C5253", x"5A564F54", x"515A5459",
									 -- x"584B5351", x"4A484F4E", x"47494343", x"484A493B", x"434B5251", x"4F565D5A", x"51514459", x"55544D50",
									 -- x"4F55515C", x"5A5C4F4D", x"5C654660", x"59515541", x"534D5456", x"4B4B5045", x"5B616057", x"70545C71",
									 -- x"566A6980", x"606DB8C2", x"6D717C74", x"5E5F503D", x"374F534F", x"4E495B48", x"5B565253", x"89715C73",
									 -- x"5B526459", x"53485869", x"64536387", x"5746594F", x"4761505F", x"704F3247", x"5E74583E", x"7C4E405D",
									 -- x"99CB8182", x"474F535C", x"435A5240", x"79754F5A", x"5F4E3D34", x"243E323F", x"474F5657", x"4D4A4C4B",
									 -- x"5B52483D", x"3B293D4B", x"54514947", x"3D404548", x"41333842", x"48535C49", x"5A4D5D4D", x"3750574F",
									 -- x"3C4A5153", x"50634240", x"50594F4A", x"55544C51", x"3B607C66", x"60605F58", x"5661544B", x"273B3B41",
									 -- x"3B214952", x"3E323E29", x"493F3436", x"18323216", x"2D44464C", x"50504F4B", x"5E5A616B", x"7B6E835C",
									 -- x"4E3F4047", x"44464B46", x"3E3E444C", x"48444B46", x"4B43404D", x"4C4B403A", x"3032333D", x"453C3746",
									 -- x"4546484A", x"4B494A51", x"4F5C4F4E", x"52534C5D", x"615E5C56", x"51505B53", x"4C483128", x"3D4E5055",
									 -- x"5054534D", x"4A4F575B", x"54525953", x"504E4740", x"4140474F", x"45494D4C", x"5C565858", x"5458524F",
									 -- x"4E605F4F", x"52554D52", x"56596061", x"5955595B", x"625F6160", x"615A5B5C", x"585B5D59", x"585C5C5A",
									 -- x"5B56555A", x"5E5C5551", x"54555256", x"54505456", x"504A4B4E", x"4B494A49", x"43383F36", x"3B41354B",
									 -- x"30383F42", x"4840493C", x"38424743", x"41414348", x"3915374B", x"444C442B", x"2A211D17", x"15151C1D",
									 -- x"08063141", x"4449423D", x"45403D44", x"3844353E", x"3731293F", x"3B3B3438", x"37364447", x"44414246",
									 -- x"4A444546", x"5549423E", x"53524B53", x"3E394042", x"4B474C3E", x"3E333F58", x"45534168", x"5E3B6267",
									 -- x"5D4B5550", x"5F625351", x"665F6A5C", x"545F624D", x"42414B4A", x"48454255", x"552F394C", x"3D404A42",
									 -- x"474B4046", x"3D3D3542", x"392D2D3E", x"3C3D3B3E", x"4B4B4344", x"45464249", x"47442A37", x"3F423C3E",
									 -- x"404C3C45", x"383F3D40", x"393F4E44", x"4B384643", x"33383C3B", x"3C3E4947", x"4463442B", x"364D3A35",
									 -- x"3A433D44", x"433C4244", x"4E494641", x"474E4235", x"4152454D", x"5746454F", x"4143474D", x"55555C69",
									 -- x"52506F5B", x"54445A48", x"5357564F", x"51565E56", x"494A5153", x"4B484E56", x"554C514E", x"483E4D5E",
									 -- x"3E52514C", x"4340372D", x"4C3E4144", x"54593246", x"5F51504A", x"4F4C5D52", x"3E3E3534", x"41444439",
									 -- x"514F4B44", x"4862755A", x"5862464F", x"5855504E", x"55695968", x"6775866A", x"615A6D77", x"56395C65",
									 -- x"6766657E", x"71676F73", x"8F6F5E5E", x"574E4A6A", x"66556B5C", x"53619C78", x"59737455", x"78605174",
									 -- x"8CA25659", x"54685A55", x"51585F49", x"568C5841", x"4246485B", x"5151493B", x"594C3921", x"3E42392E",
									 -- x"3D473747", x"4449474D", x"3540483C", x"4C443D3D", x"4B40414E", x"4E567953", x"4F505851", x"4F596852",
									 -- x"365B5D4C", x"60714B4F", x"55464945", x"405B5856", x"63726955", x"4D574E56", x"58655554", x"5656363D",
									 -- x"48323744", x"57553A51", x"5A90705A", x"434D595B", x"596B4F4F", x"414A5C69", x"61646662", x"6F58525A",
									 -- x"53453E3E", x"3C404440", x"3B404946", x"483F4840", x"40454B4C", x"3F484941", x"4245484C", x"4A454C5F",
									 -- x"4C4E5455", x"4F505554", x"57605D5A", x"5D5A575F", x"605F5247", x"52535B55", x"52423E43", x"4853564A",
									 -- x"5258564D", x"4A525A5C", x"53514F4C", x"49463530", x"2B375456", x"4D54645A", x"62545757", x"5A5E6060",
									 -- x"58646156", x"5F64585B", x"61606464", x"5E5B5E5F", x"635F5E56", x"59565956", x"5E5C6057", x"53575255",
									 -- x"59585655", x"55544F4A", x"524D474D", x"524F504D", x"47474B4E", x"4C4A4844", x"44364A4F", x"47342E65",
									 -- x"92324F5C", x"49513E42", x"3D3F4444", x"3F3F4345", x"2A393C52", x"52443F2E", x"23181115", x"171F1B0F",
									 -- x"00131820", x"48483732", x"33323D3C", x"2C362F35", x"36435148", x"3D464A45", x"58494B56", x"54555764",
									 -- x"5D62585A", x"473D3445", x"3B4C3946", x"5D4F4048", x"6B4D595F", x"543E4880", x"6B534A71", x"689D7A95",
									 -- x"77655235", x"737E6686", x"7F759D6E", x"7C758160", x"58514D51", x"665B476D", x"45251432", x"52544E4C",
									 -- x"4A4A374D", x"4D474D47", x"45474340", x"3C48473F", x"3E3D3E52", x"59594A45", x"3E3F3C45", x"4C4A403C",
									 -- x"3F3A2D39", x"393F3736", x"2C333F32", x"3826322D", x"383E3731", x"38413E49", x"393B324E", x"4140433D",
									 -- x"4947414B", x"433E4C50", x"473F4E4F", x"464C473A", x"3D453933", x"45383749", x"404C5D50", x"5C474B47",
									 -- x"504E6250", x"4A3A534E", x"5458584B", x"54525356", x"594B4E59", x"51434857", x"58525C51", x"4F49516E",
									 -- x"5A565448", x"4E3A505C", x"50494A45", x"62504E54", x"4B504D59", x"4A45403C", x"393F3748", x"4A46414F",
									 -- x"4445404B", x"4C3F4A4E", x"5B3E4D50", x"414A515E", x"5993595F", x"60534C57", x"4C472C6F", x"46245952",
									 -- x"5660A099", x"6F7B516C", x"80595255", x"5F5B5667", x"734E4E59", x"716F715D", x"686F4F5B", x"5741434B",
									 -- x"404E615F", x"6F59666B", x"57495B60", x"275A4E35", x"4A404645", x"45445039", x"45494B39", x"5048475D",
									 -- x"4745432D", x"74323B48", x"43394538", x"4A5D4A53", x"4962556F", x"595C5062", x"5A563F40", x"47586345",
									 -- x"43405A5B", x"5F485959", x"4949555B", x"3D56646F", x"5D6F5F4E", x"47575446", x"5C605D58", x"7E603A3F",
									 -- x"4C6B575C", x"9F979E63", x"779472A0", x"916AA49C", x"545D5552", x"4B425B76", x"7F4F4D4D", x"57554542",
									 -- x"4B433F3E", x"3D40423D", x"43454B41", x"4C47544B", x"4D585351", x"4E514E56", x"54585650", x"4F535451",
									 -- x"58555956", x"4E53564A", x"5B595E58", x"59575F60", x"686D6E65", x"65687159", x"5357646D", x"69615A54",
									 -- x"5C646358", x"53585C59", x"605C5358", x"616F6870", x"575E7864", x"55505836", x"534A5B62", x"6762605B",
									 -- x"50525D5A", x"545B5F5F", x"645A5657", x"56555450", x"4D4F534D", x"5555564C", x"4C414B48", x"47484353",
									 -- x"454A4C48", x"494D4E4B", x"4C4A4549", x"49454B4E", x"504E4F4E", x"4B4C4E4A", x"4B4E453F", x"4D4F3D35",
									 -- x"404A4849", x"3D3B3B41", x"453F4144", x"40404544", x"4E4B504D", x"393E3225", x"1C1E331D", x"1803120A",
									 -- x"05150C24", x"50464847", x"4E567559", x"50505143", x"67576D54", x"5F566255", x"49484953", x"49514444",
									 -- x"4B484F63", x"1D313937", x"182E5027", x"1E2E0D18", x"1A2B4325", x"1B3B3C43", x"4F476A5C", x"6983767B",
									 -- x"59626B57", x"7A5E4553", x"4E5C6442", x"5F503E66", x"5C435B65", x"51444F78", x"3730321A", x"58304850",
									 -- x"473B306E", x"79586550", x"6C7E6F5F", x"5C5B515A", x"4A535255", x"56665E4F", x"4E475345", x"57505855",
									 -- x"5553554B", x"4D494D4A", x"4B4B4A53", x"50433F3D", x"443D4444", x"37464341", x"4245393F", x"48444847",
									 -- x"3D444632", x"42484048", x"514C4841", x"494D3F40", x"4C4C364D", x"4D486958", x"76725D4E", x"4B444143",
									 -- x"54494550", x"4E424144", x"524C3F36", x"5555474C", x"554A494E", x"4A43464C", x"51624F5A", x"4B703F4C",
									 -- x"595F564D", x"504D5D5E", x"534F484E", x"5550604B", x"3D554B46", x"2E384041", x"4D3B3C57", x"483A3B3D",
									 -- x"3E534E36", x"30544752", x"4640484B", x"3D283E4D", x"4D535B49", x"43423A4A", x"45466061", x"484A3F53",
									 -- x"52516070", x"64645A52", x"644F4E5A", x"615D7B86", x"5B5A6562", x"65645254", x"5F7B6549", x"5151444C",
									 -- x"64586567", x"5859514A", x"4B3C375C", x"6B5A5D56", x"85606F4A", x"4E4C5032", x"3A2A3845", x"4E5C5859",
									 -- x"695A605E", x"4E405E4C", x"68434F46", x"31614250", x"512B3931", x"4D554649", x"3348606E", x"34454A27",
									 -- x"22364852", x"4D2F4C55", x"47574762", x"50555D5C", x"675C4949", x"4E475E55", x"5D535438", x"2B303734",
									 -- x"334F3835", x"311E412D", x"23152832", x"3520161F", x"2D2F3E25", x"36233D4A", x"4F3A404E", x"4F477271",
									 -- x"494C4849", x"434E4943", x"4F565C50", x"575C6057", x"5A535D57", x"56535858", x"59624F51", x"594E5256",
									 -- x"5C575349", x"55554E4F", x"6B5B5756", x"54556464", x"6964625C", x"55565559", x"5A504C5C", x"5C5E5F6B",
									 -- x"6A646567", x"5C636269", x"7A595663", x"6C5F6060", x"44515361", x"576C4B53", x"62736462", x"5F5E675A",
									 -- x"59615557", x"575A5D56", x"59564B4F", x"4D444846", x"4F544647", x"4E494B47", x"3B403D3D", x"433A4546",
									 -- x"453E4251", x"473F534E", x"46574B46", x"42464C4F", x"42465D42", x"4C504244", x"5346463C", x"3F453633",
									 -- x"27343325", x"3A36343D", x"46443634", x"4A4C3E4F", x"494C514A", x"452C1B11", x"131D221B", x"1A081717",
									 -- x"13232C39", x"68554C67", x"6A637E5E", x"5B5E493C", x"47444547", x"4D3E5049", x"3640243D", x"332B3A41",
									 -- x"380C1553", x"1C3B3630", x"3829354F", x"4330353A", x"3E52452F", x"28363F2C", x"3E463047", x"53384C43",
									 -- x"414F7B68", x"3A41412A", x"32423751", x"4D3F4D53", x"5E536650", x"3D483D2F", x"575E5839", x"18232835",
									 -- x"631B495E", x"594F4543", x"4D747367", x"49636C51", x"45464958", x"574B5950", x"4E53505C", x"5754545C",
									 -- x"5955645C", x"5E535F57", x"5A63565F", x"64665E57", x"535D5A59", x"52564D47", x"46523F45", x"4D504743",
									 -- x"44304545", x"38444B4B", x"4C363E4E", x"47473E42", x"534E4648", x"5859554B", x"3D384043", x"3D3D4450",
									 -- x"4A49393A", x"4A41353E", x"5A4C433F", x"52494D51", x"3A324349", x"3E3F484D", x"505B5B52", x"515B494B",
									 -- x"56392266", x"593B5E47", x"53324A5B", x"4A43363D", x"2A484244", x"503A4857", x"48474545", x"413A3C42",
									 -- x"40393C35", x"4C534948", x"4E473141", x"49584665", x"50444E4A", x"443E4241", x"48423648", x"3A454C48",
									 -- x"4F4D3D57", x"48494D4D", x"51473A53", x"55515956", x"666A745C", x"5A5E606F", x"5943546C", x"6C55627F",
									 -- x"686A5953", x"4A524F55", x"604A4E5E", x"5F536156", x"554C5750", x"5063594B", x"624B434C", x"455C4B47",
									 -- x"4C455952", x"50303F4B", x"58373E5A", x"5348424A", x"462D3A43", x"345C6C52", x"4D34515A", x"4A713646",
									 -- x"63694641", x"52574F51", x"525E4F57", x"6367635F", x"46585A60", x"5044535C", x"5C384D44", x"3A3C4F44",
									 -- x"55595453", x"5937403C", x"40294D5A", x"2423383D", x"544C5151", x"3F614544", x"515E595E", x"34495B5B",
									 -- x"54505053", x"56525457", x"5E595A55", x"57515557", x"414E4F4B", x"53505B5B", x"60776363", x"615F5A66",
									 -- x"665F5B52", x"41535D57", x"575C665A", x"71585D53", x"575D5156", x"4C59544C", x"59534553", x"59676470",
									 -- x"6A695F62", x"66646264", x"625D615F", x"59586060", x"71515756", x"38606266", x"786F5659", x"58575F5D",
									 -- x"56646259", x"4F4C444D", x"4C434941", x"4E494F4A", x"444B4743", x"42424541", x"37404137", x"3E363F38",
									 -- x"363C4F47", x"3D42454F", x"4C40433E", x"4D4F403A", x"36404A3A", x"3B343D4B", x"3A2C363C", x"2D464137",
									 -- x"4526444D", x"4549484C", x"4540464A", x"3F4B5A4A", x"53554E62", x"5F582E19", x"24282243", x"25413C3A",
									 -- x"40485B4D", x"4A4C5457", x"593C494F", x"544E4A3F", x"4A484445", x"3A433D41", x"2C204049", x"40406135",
									 -- x"413F3D4C", x"42360E3F", x"3F3A4250", x"46455D4F", x"432B2B35", x"1C3E4830", x"35333C36", x"1B312C3D",
									 -- x"371D2B3B", x"422E3937", x"383F4633", x"3A273734", x"32372D24", x"3835244C", x"31363D3E", x"4A5E4060",
									 -- x"544B6052", x"3B3F474D", x"363A494F", x"4946402D", x"4F524839", x"4A52444B", x"56484155", x"5D544E4D",
									 -- x"4F483E41", x"3B394943", x"4C545058", x"4F4F5456", x"566A6D5B", x"5A5F5852", x"6B55474D", x"606D6354",
									 -- x"654F6271", x"65526454", x"686B5E51", x"6D795C61", x"584F4C68", x"5B65584E", x"38455442", x"44433E44",
									 -- x"4B34473F", x"453A4650", x"4547484F", x"524E4248", x"45505C69", x"5E56535A", x"5F57585D", x"48576255",
									 -- x"5086604E", x"543A4D60", x"524D514A", x"4F4A5364", x"4F4C4757", x"4D595760", x"4E515E47", x"38414441",
									 -- x"494A464E", x"4C49494A", x"3F412336", x"44454446", x"5F494447", x"46474E46", x"3A675636", x"2F493D44",
									 -- x"4651474A", x"4F41403F", x"4B47424D", x"4756413F", x"55525344", x"555E565D", x"614B5B5A", x"5062585B",
									 -- x"45585554", x"45434259", x"5759535D", x"2A5B5C33", x"2D495741", x"46382E4B", x"5B49384D", x"56435552",
									 -- x"52523A44", x"4B3F3243", x"41372B44", x"4B3D3D43", x"426C3750", x"3E3A3C40", x"4C623C2E", x"5A624C4A",
									 -- x"59502F2D", x"435D555E", x"524D6070", x"5D606E62", x"617E7756", x"63616152", x"484C4245", x"42294147",
									 -- x"524D5640", x"444C3F3F", x"5349314A", x"513F424E", x"6544474F", x"4F4F504F", x"65715B52", x"525A595A",
									 -- x"615A5B58", x"60575D66", x"5B60655B", x"57545C5E", x"5E7A6F66", x"6B5F635C", x"66647D79", x"6D6E7D66",
									 -- x"615F4E3B", x"2D4F5664", x"56665769", x"5E615456", x"5C60616B", x"645C5F5C", x"6A6B5952", x"5B615B61",
									 -- x"565D5758", x"58575F56", x"4D585D58", x"4D545650", x"464B4D52", x"4C575546", x"51555554", x"46454445",
									 -- x"4336414F", x"29474C4F", x"44384337", x"4144423D", x"2D314045", x"43474642", x"3B484440", x"35313439",
									 -- x"2E3E3744", x"433B4539", x"3E513544", x"3C47393F", x"4046473B", x"3E203E48", x"30294143", x"4C464647",
									 -- x"4B4F5064", x"4B436262", x"4F5E5E5A", x"54576963", x"5A5F576F", x"6D73564E", x"4B5C635A", x"594D4756",
									 -- x"58665C5E", x"5B546555", x"56495163", x"55496060", x"4A464F4D", x"5B5D6564", x"576C7884", x"5F655C60",
									 -- x"5E4A5461", x"5848415B", x"614C4C3F", x"47515445", x"554B5862", x"47463B44", x"413F4128", x"202A373A",
									 -- x"37383D31", x"3D3D4A52", x"3D484D5E", x"464B2E38", x"2B343A37", x"32354D80", x"2C454255", x"647F6957",
									 -- x"5D57413C", x"51514B43", x"4A3F4543", x"4143423C", x"3B414F34", x"5A555355", x"3B484D46", x"4348534A",
									 -- x"455D4D4A", x"43494046", x"4C46444F", x"47444644", x"42404942", x"4C444455", x"4D614B33", x"4F624A59",
									 -- x"5A576A4C", x"615D5568", x"4B5C6C59", x"5F725E5C", x"5B5A6560", x"59525A58", x"5B5C4E52", x"50365B3E",
									 -- x"414D484C", x"4B4E5A3A", x"4C4E5C54", x"57514D55", x"4C524843", x"5159595A", x"66534C56", x"50465E62",
									 -- x"5D4B5938", x"49665255", x"59655459", x"56564E56", x"4D4B3E4A", x"4250434F", x"4F4C5559", x"58596754",
									 -- x"43585448", x"464A4640", x"4C4F4E4C", x"4D4F494D", x"46484848", x"3B475338", x"4F4E4D43", x"4D5B5357",
									 -- x"50685E73", x"605E4F53", x"504F585A", x"444A4655", x"634D5050", x"57534845", x"414A4A5B", x"695B2A55",
									 -- x"46444741", x"594A4748", x"5B675A68", x"5D635069", x"57676F59", x"6D4F3B4D", x"4C445C60", x"5B525B5F",
									 -- x"563E4F5B", x"484A654F", x"3E47313E", x"42404D3A", x"3E2C4B4B", x"5C4A3F39", x"4B2D4452", x"5D5D5B42",
									 -- x"35434A49", x"495F5E77", x"5B535F5C", x"4D54615F", x"5D504A41", x"65655C50", x"5E736356", x"5341443E",
									 -- x"4A443F4E", x"51565D61", x"6C5C505A", x"61615252", x"45615541", x"5549525F", x"55696459", x"68615E5E",
									 -- x"5E5F6469", x"77746E69", x"5E686E69", x"68696A67", x"5E736B64", x"67646864", x"6D676E59", x"5F5B6159",
									 -- x"57634E56", x"585E6664", x"64595862", x"595A6962", x"5E5E6169", x"64636870", x"606E684F", x"5A514E52",
									 -- x"5351504F", x"45535B4B", x"4D525050", x"45453D39", x"3E484B35", x"40402E47", x"42404645", x"3E453F3F",
									 -- x"3F45515F", x"54554344", x"3B35383A", x"333A3434", x"32293E48", x"43433E3B", x"3B41413E", x"4443433E",
									 -- x"542C2A3E", x"37424634", x"41433E48", x"42373F40", x"4F47463A", x"4E2C5150", x"3D4E6048", x"53585C54",
									 -- x"565B6578", x"546D8C5E", x"647C766B", x"76696474", x"58595754", x"54515359", x"54525E5A", x"52555258",
									 -- x"5D636464", x"615C5A5F", x"56534957", x"5C5A522E", x"4344304E", x"55596162", x"5A585032", x"59464C61",
									 -- x"3E4B4144", x"42475A4B", x"3F3A4843", x"534A4853", x"6257473B", x"4C403A56", x"4B52445A", x"4C51563E",
									 -- x"3B3A4434", x"33422B3D", x"4131443A", x"483C3D3E", x"2D334E31", x"4635555B", x"40555165", x"56434945",
									 -- x"45564836", x"4C454541", x"40423D43", x"3A44433F", x"3B393C4E", x"4140443C", x"49484841", x"42404D46",
									 -- x"5E46475C", x"484D444D", x"4847494D", x"42393F4C", x"473C3F32", x"3238383B", x"36253E5B", x"3E4B504A",
									 -- x"493B4F4A", x"534B556B", x"4F4A5350", x"526A5455", x"474E4D51", x"645F4F54", x"555B654D", x"4F517254",
									 -- x"49664C5F", x"66575143", x"545A5459", x"435A4D60", x"54555C4B", x"57535053", x"565B5941", x"504B5E56",
									 -- x"43355457", x"55503E3E", x"554C4C48", x"5448504A", x"4D465240", x"40493C4F", x"4339584E", x"4D534E55",
									 -- x"55414C49", x"42444946", x"43434E44", x"3A43404C", x"2F49394B", x"5A443A53", x"534C5542", x"53566160",
									 -- x"50525A69", x"56556364", x"62615057", x"724F4357", x"602E3448", x"4F4D4F47", x"4F554F5B", x"4C474047",
									 -- x"53504452", x"515E5455", x"4D384A4C", x"4648504F", x"4D385F5C", x"57516045", x"5BAB887A", x"A99F6267",
									 -- x"52535B3B", x"46464D38", x"463C2659", x"3D47514C", x"404B5950", x"5E544C4C", x"5D593D4F", x"635C5A4D",
									 -- x"535F6250", x"45556579", x"6A555051", x"5B565B7F", x"594A6067", x"63635B58", x"5F527752", x"4E6F5A5C",
									 -- x"61424C67", x"6E685862", x"66464D4D", x"39505D5F", x"616B5854", x"585D5E55", x"5A515551", x"5B616B5B",
									 -- x"62686663", x"5A5E6572", x"776D666B", x"6F6F6E72", x"6767645F", x"5D676E70", x"666B5F63", x"5F6A5E6B",
									 -- x"73526B6A", x"666A635F", x"665B6B67", x"6B6D7D68", x"77756456", x"4D61565A", x"465A5A4B", x"524E4A4F",
									 -- x"52474348", x"4B573D3B", x"4B4E4B4F", x"47443A3A", x"4B50464C", x"41283942", x"463F4F4E", x"463F435B",
									 -- x"48515247", x"56383536", x"34343446", x"3B3D4447", x"5D4C534A", x"3B434B4D", x"3E465944", x"55495249",
									 -- x"48564B49", x"4B5574B4", x"8542504D", x"525C5B62", x"76675F53", x"5F4D6059", x"5A536076", x"585A5A61",
									 -- x"6E4A7152", x"38826A68", x"6365786B", x"6B645758", x"534D504A", x"5C575F5F", x"5A555454", x"4F5D5760",
									 -- x"50554252", x"504B614C", x"4E5B5046", x"4B50514F", x"56472F4F", x"564F4C57", x"4E434143", x"39414E46",
									 -- x"4D5D485A", x"513F4959", x"69514E50", x"583F3F3E", x"45393036", x"4D46453A", x"47434D4C", x"2F3F413B",
									 -- x"3B333D3B", x"3740222C", x"32332A29", x"263C4643", x"47383633", x"343C3F2F", x"253D4331", x"3F3D3E4D",
									 -- x"4C464247", x"442A2947", x"49432F42", x"3D313A38", x"51363545", x"3138453A", x"49484541", x"4B4D5347",
									 -- x"394A4144", x"3E4A4C47", x"4A494744", x"433A3E52", x"5A494E4E", x"3B424039", x"40393C45", x"352E424E",
									 -- x"3D384B34", x"3250474E", x"54344A5D", x"38504C43", x"3E35453E", x"69514A4D", x"4C515132", x"49464A4D",
									 -- x"37485249", x"605D596F", x"605D625E", x"5D656265", x"64526363", x"6767555E", x"62515A59", x"5C4F5057",
									 -- x"54585C5F", x"5B5C565A", x"5F5E555A", x"53625F6D", x"5C5F585C", x"574A765D", x"4C554734", x"46544D35",
									 -- x"444D3B3A", x"4547434C", x"3A392837", x"333A4440", x"3D3A2C4A", x"54494B54", x"483A4B40", x"2C3E6543",
									 -- x"47545C76", x"626E655E", x"5C4D3F3F", x"4F414755", x"6249515D", x"5F524E4B", x"534B5454", x"39435638",
									 -- x"47484D58", x"4A595950", x"46483D2F", x"3E514546", x"544A4E3F", x"58595842", x"597C5C46", x"5F876155",
									 -- x"5D43575F", x"3C454F60", x"5B4A543D", x"4A47684D", x"45785A50", x"49595145", x"4C575263", x"5A565660",
									 -- x"576B7367", x"62647573", x"63615645", x"44404670", x"674E6061", x"61636061", x"66605B51", x"433E5B49",
									 -- x"604B4F65", x"7468533F", x"4F484C6D", x"61525A56", x"4E5B6164", x"5A685E50", x"5C546763", x"4F566B61",
									 -- x"57555864", x"554F4A4E", x"4B535A62", x"5E5B5350", x"584E4E4D", x"454D4E52", x"55585968", x"5D5C5559",
									 -- x"462C5E60", x"6D665857", x"59665C63", x"537E635B", x"61606046", x"574D4F54", x"58605757", x"4D504548",
									 -- x"3C404955", x"67592438", x"464B494C", x"4D463226", x"443B404B", x"4755564E", x"4A3D4544", x"584F4545",
									 -- x"3E402938", x"454E5156", x"46414657", x"544B5D5B", x"474F6360", x"535E655A", x"57525659", x"594F4F61",
									 -- x"59675D6E", x"5C58645B", x"6C5D5E5C", x"6E755A5C", x"5B5B5960", x"5D63635E", x"54515868", x"514B4951",
									 -- x"54554E51", x"4A595058", x"524C6854", x"5159514B", x"5A545253", x"605B554E", x"5558573C", x"56403B42",
									 -- x"493A343C", x"52564F4E", x"444E4F4F", x"5C4F495E", x"4D314147", x"5C4C3649", x"363A3B4C", x"61503C3F",
									 -- x"3A4A4941", x"34454544", x"4D2C554C", x"3F4A5060", x"4548444D", x"46454936", x"32383F2F", x"56583E32",
									 -- x"3B464237", x"36373F36", x"36424349", x"42414736", x"45454A5A", x"1E2C375B", x"4E4D4734", x"423B4841",
									 -- x"4F423941", x"41503B35", x"26313346", x"4E2C3C32", x"4129462D", x"3B3D4744", x"1E36392E", x"31363A31",
									 -- x"2D392C46", x"3B395C41", x"4C484842", x"463D3538", x"4336445F", x"4A444745", x"4D5C614F", x"5B4B5D55",
									 -- x"4A5A3242", x"48414047", x"473A3447", x"444D3131", x"4043494E", x"3E544A4C", x"40393D49", x"5240495A",
									 -- x"5B574F48", x"46535446", x"4E51475E", x"52665956", x"48434F60", x"657E5B55", x"5F635D5E", x"5B5F4552",
									 -- x"54505247", x"3A5F737E", x"63768378", x"8B79605D", x"6574556F", x"71598461", x"53606744", x"4B664C50",
									 -- x"2B624347", x"4A534C42", x"47403748", x"45483F3A", x"4E4D3B3D", x"454B4B40", x"2E342737", x"3C47483C",
									 -- x"464D4D2F", x"4F45483C", x"48444C49", x"475F443C", x"43525450", x"6155484A", x"47455047", x"524C4E66",
									 -- x"5A444C36", x"3F43604D", x"50494249", x"4E443C51", x"3C374138", x"37465B50", x"4D424C2F", x"3E55323C",
									 -- x"6E4B4C61", x"525D4F57", x"55555954", x"5C543F3A", x"57445148", x"435D543E", x"5F4E3C52", x"5B5B5B4F",
									 -- x"5A7A8C8A", x"7D67695D", x"6D775C5D", x"7F815A61", x"54516347", x"59505D73", x"65645852", x"54555D56",
									 -- x"52584C61", x"6A5B6B59", x"5A56545F", x"55504E50", x"444A554D", x"5D6A5D5A", x"5C52595D", x"5B635F52",
									 -- x"4C363444", x"4B504937", x"3A494840", x"38495357", x"50544F54", x"5256585D", x"5B665D5B", x"74626674",
									 -- x"6269585F", x"74547A62", x"65656361", x"5785645C", x"5E6A6C62", x"78444B56", x"685B5759", x"4D474542",
									 -- x"4745422D", x"3B363252", x"474A4947", x"4C3F2D22", x"2F433558", x"5C6A6950", x"4A4C5544", x"6054534F",
									 -- x"0E2F103D", x"59713E4C", x"64575C66", x"615F665E", x"5C5F6464", x"606D807B", x"755D5370", x"787B6776",
									 -- x"6063625F", x"576E5D54", x"4D6C624D", x"6E575E58", x"4E575962", x"5758564C", x"52414147", x"4A29314B",
									 -- x"44293447", x"3F4F494B", x"4A50624A", x"504F4D56", x"4A4D4F52", x"57544F50", x"574E4D4D", x"55525549",
									 -- x"4C524B4C", x"5D494B52", x"4D4F4D49", x"533F4258", x"51485D5E", x"5B5E3651", x"4A324A56", x"44373946",
									 -- x"383B392D", x"4A4A4045", x"36214A44", x"414F393E", x"3B43403D", x"3B3B3938", x"325B463E", x"483A3240",
									 -- x"4E533C3D", x"453F4742", x"41434A52", x"4D3E402A", x"413C433A", x"473F3751", x"56625E44", x"373A5C39",
									 -- x"413C474B", x"44414143", x"50625E51", x"513D5145", x"44455847", x"45513F41", x"393E3134", x"372A232C",
									 -- x"2F461F27", x"39444F3D", x"3C3D5249", x"3C363630", x"2C39424F", x"48464C3B", x"4A363941", x"5A505958",
									 -- x"545E585F", x"58655053", x"594E4B55", x"4E4D4F52", x"4E46514C", x"49605B4D", x"4D48766E", x"4759565D",
									 -- x"6F5D3F66", x"4F53603C", x"47433B4B", x"52555C4E", x"4E5D5852", x"4E5D5B64", x"5F604F5B", x"635C4861",
									 -- x"5565534E", x"565D6864", x"66736060", x"64625962", x"574F5150", x"554D4254", x"5858555A", x"5C624F57",
									 -- x"4D495D73", x"5454634D", x"5E56625E", x"5958474E", x"684C5056", x"47455143", x"3E434349", x"47534D3B",
									 -- x"404F4435", x"44423439", x"405F563B", x"39442046", x"4A4B3B30", x"494E4B47", x"313B544E", x"5548444D",
									 -- x"52545A57", x"5253544B", x"4F4C5252", x"482F343D", x"463E343D", x"424D5050", x"4A3F3639", x"5E4A424A",
									 -- x"3A505437", x"4248462C", x"42473F2F", x"444E3E38", x"5F474552", x"41444356", x"6D54614E", x"4A684D41",
									 -- x"6D6B5F63", x"60635F64", x"5C716580", x"88693F58", x"505E6B46", x"625B554A", x"5A694D5F", x"69716D64",
									 -- x"66616761", x"575C5B76", x"60595C49", x"39525358", x"5533494B", x"42385067", x"635B625D", x"5B63686B",
									 -- x"4E4E615C", x"50515F52", x"5055545C", x"5D6A6B6C", x"68765D5D", x"5A575D65", x"645F535E", x"5E565D51",
									 -- x"68545347", x"5055795D", x"6248636B", x"62856857", x"587D5C73", x"714F464E", x"4C324444", x"4B3B514C",
									 -- x"4C4F6449", x"4B455142", x"45484E4C", x"53495363", x"53584C70", x"55565862", x"60606A63", x"8B6E6C6B",
									 -- x"383F3B54", x"667A5655", x"7462626F", x"6071645D", x"72655C63", x"5E555B53", x"5251685F", x"73645B52",
									 -- x"4F66514D", x"454E4E4C", x"4C48424F", x"46434B49", x"4C50514D", x"4C3E4F3F", x"423C4B5A", x"4B3C3E38",
									 -- x"28413F5A", x"55454A42", x"454D5E51", x"4F393D4A", x"3C414945", x"493C3B3C", x"34463731", x"37354256",
									 -- x"5952604A", x"474D513B", x"363F4039", x"463D4D4E", x"46495D42", x"47403647", x"5341403A", x"3944283E",
									 -- x"50454742", x"66444635", x"3E59444C", x"52383835", x"3230412E", x"302C3D4C", x"3334423F", x"3920433F",
									 -- x"3A524345", x"47503B3C", x"34393F49", x"4F605F43", x"47434D3F", x"27484B54", x"543C3C35", x"3B38373C",
									 -- x"3F44573B", x"3A253E34", x"3D4D443D", x"3E42473D", x"47434845", x"4A514E41", x"45513B33", x"3535303C",
									 -- x"32464047", x"44403450", x"35294441", x"36424D39", x"393F3A49", x"55414942", x"5A4C5057", x"49473A3F",
									 -- x"44514C46", x"5359346D", x"6B564F5C", x"6C5E5E52", x"6D56504D", x"4D52526D", x"65584F4D", x"2F4C5952",
									 -- x"4548505D", x"4B567556", x"4D4A3951", x"52586255", x"5A665E5A", x"64404C61", x"58535052", x"5B617568",
									 -- x"56587056", x"555F5153", x"51545361", x"58445A5F", x"5D514D54", x"462B4A5A", x"53485765", x"58615373",
									 -- x"5E476E57", x"5C595A65", x"595C564E", x"5047575B", x"5C52544C", x"52575A55", x"6E585D50", x"5C55524D",
									 -- x"484F4F57", x"51514C62", x"614F4443", x"34353B4A", x"49454D4B", x"413F5556", x"58544D52", x"56475651",
									 -- x"5E5C5752", x"5F5B5757", x"5662534F", x"48403F40", x"57534558", x"4D473E4C", x"4F39505A", x"67555156",
									 -- x"4F58574C", x"55394837", x"44353843", x"5652453D", x"48414C5A", x"463D4059", x"4F4B4259", x"555D6067",
									 -- x"6C573F4B", x"4A59485B", x"60695A60", x"44555C5A", x"62586667", x"6F5D5F67", x"5D603E61", x"52554E56",
									 -- x"636A5D59", x"4649404F", x"656F5D55", x"4D535D5D", x"514A525D", x"6F635B64", x"604F5D58", x"555B615A",
									 -- x"566C655E", x"6D675C6A", x"64646D64", x"63605D54", x"52544C53", x"56475065", x"53504F51", x"584B4F50",
									 -- x"60636254", x"53657066", x"5D3D706A", x"596B5752", x"536C4178", x"6C553B65", x"4F54565A", x"675D6153",
									 -- x"5A434238", x"46545147", x"54534F41", x"5F5A5460", x"58435F60", x"4F3E5A64", x"73666D66", x"4B3E5758",
									 -- x"5F606A5A", x"6D6F6958", x"575D5050", x"5653544F", x"4E4F534D", x"4F3E353B", x"51454E4C", x"30393837",
									 -- x"413A433C", x"453D424B", x"453E3C43", x"47434144", x"47594337", x"3B4F5E38", x"426C7A57", x"3F494B40",
									 -- x"45514B42", x"49494243", x"4348353E", x"4D5A3758", x"3B3E4836", x"41393537", x"2C393C30", x"1F36473F",
									 -- x"40413E2E", x"2D33423D", x"35351F2E", x"32232941", x"381E2B49", x"291F3030", x"34313B2D", x"2F2B2A38",
									 -- x"393D4B4E", x"44323A35", x"3D472241", x"3237383D", x"39372D2A", x"1A303330", x"2C2C3B42", x"4D383C32",
									 -- x"3B414246", x"4B454048", x"3839484C", x"4F4F5A8B", x"52444D52", x"534F5D5E", x"403E4533", x"353B3D3C",
									 -- x"3F4F483F", x"37363B2C", x"3A3F3C3A", x"2E3A3E3E", x"21464738", x"49393E2E", x"483C393C", x"26504C36",
									 -- x"2F5A5532", x"353E3643", x"3C4B3B3C", x"43463736", x"42353A3E", x"3C4E4340", x"3D473946", x"4F514532",
									 -- x"5255473F", x"404B5566", x"523E474E", x"4A4B4A4F", x"4C4A6453", x"4D3A4C44", x"573C4432", x"49484E53",
									 -- x"493F3C41", x"3D565954", x"4D4B434E", x"50526057", x"50575C50", x"47554E5D", x"5D4F4B59", x"52515656",
									 -- x"5C42525A", x"4B493F53", x"3D495958", x"533B5365", x"534E5259", x"554F5A58", x"4C595A70", x"6058535C",
									 -- x"4F494A46", x"4B524746", x"4053323D", x"414C5557", x"52575957", x"6F765F63", x"6D5D6553", x"575C5E6D",
									 -- x"76635970", x"4E616262", x"645A5C60", x"44484F4C", x"5E38575A", x"474C5552", x"615C6052", x"586F656E",
									 -- x"68606354", x"5F5C676E", x"5F5E6D67", x"66676A79", x"5F585F68", x"5E5E525E", x"51667B68", x"6A667264",
									 -- x"6D65617A", x"675D6D5F", x"64646657", x"6B465053", x"59505050", x"39533D42", x"4F676861", x"515C615C",
									 -- x"725F504C", x"51686164", x"7750625B", x"4B534C63", x"5B61505C", x"59394770", x"5D2E554E", x"5846595A",
									 -- x"5E5C5257", x"4D5C4F4B", x"475A4B53", x"4E51525F", x"65575E5B", x"6B625057", x"5E43585A", x"5E6D5857",
									 -- x"4E52575D", x"61615A52", x"57575D51", x"535F5A52", x"4F4A3850", x"414A4D46", x"4C50555E", x"51434B54",
									 -- x"49665F5A", x"59717582", x"733E615B", x"635A5E4E", x"76424D66", x"4A274677", x"59734F59", x"64665256",
									 -- x"53553841", x"5558656A", x"626E746A", x"63706568", x"5F656E69", x"62707263", x"575E6A5D", x"57705963",
									 -- x"59564B53", x"5250453B", x"55573A4E", x"43554040", x"513F3F4D", x"402F3944", x"3C403E45", x"3E5B8352",
									 -- x"40152B4D", x"3E544C51", x"58504D50", x"38404645", x"48304141", x"3E3F464B", x"61543A3E", x"484B4641",
									 -- x"3F45433C", x"41494539", x"303B2E37", x"40433A3E", x"40343A3F", x"3F4C3334", x"33263C3C", x"2E3A4744",
									 -- x"41333333", x"314E495A", x"46283448", x"38313F4F", x"40392E33", x"363F4133", x"2F343332", x"343B3143",
									 -- x"2A39413A", x"34373822", x"4F5C4B2E", x"3038493C", x"41363E2E", x"3C4A362F", x"2F374534", x"45453131",
									 -- x"40474643", x"45433E41", x"483A4140", x"40454048", x"46484E46", x"4044504F", x"43394143", x"43434246",
									 -- x"633F5B36", x"28323945", x"3D2A4250", x"35364A3F", x"363C4338", x"2F2F5D5A", x"3F483C36", x"3C3B2F4E",
									 -- x"422C2334", x"35433C3E", x"53483E46", x"43433D43", x"43393D46", x"3E3F3C31", x"41394231", x"432E4D44",
									 -- x"4149363E", x"494F534B", x"46464749", x"4A4D4A3A", x"39464241", x"42414655", x"4A4D4C4A", x"4950495A",
									 -- x"47535744", x"4750306B", x"4D426156", x"505A5C46", x"54495B59", x"655E5556", x"5862565D", x"6050565B",
									 -- x"56456F44", x"37455165", x"5E5A5B67", x"5F714D6C", x"5F636B71", x"6A8E656A", x"58476254", x"444E4156",
									 -- x"333D4646", x"403E3C47", x"724C2757", x"4D474F50", x"4F3C4549", x"3D3E5048", x"3F373420", x"46655150",
									 -- x"5C4A554E", x"575C665D", x"545F615C", x"61525164", x"65656D69", x"67656068", x"667C7266", x"6564847B",
									 -- x"706F7681", x"9267779F", x"96906C85", x"6A6E8175", x"7B727E5E", x"67846858", x"5F738F7A", x"5460565D",
									 -- x"63667441", x"595C5E5C", x"56584F4C", x"795E6173", x"58676675", x"616C7067", x"7B8C7363", x"69715F68",
									 -- x"676D5C5E", x"6E736E8F", x"57595063", x"6E515C5A", x"5F5F5D58", x"6A645A63", x"6D717F86", x"626B6A62",
									 -- x"6453645B", x"6B7A585A", x"55455950", x"5B52575B", x"59625E67", x"564E5A5B", x"5D5F5D5C", x"69614E61",
									 -- x"49555752", x"504D4D57", x"514B5250", x"53625759", x"5854505C", x"4E485651", x"4E5A5055", x"5149424E",
									 -- x"57774F50", x"5F7D8463", x"4658635E", x"574C586D", x"643C4759", x"514C7156", x"615F5360", x"4E5E4976",
									 -- x"616F6077", x"7B6D6A6D", x"70647869", x"7577786E", x"70655665", x"7567535E", x"4D5A5758", x"57665360",
									 -- x"685F4C43", x"49485343", x"744B4444", x"40474428", x"3A414550", x"5C4A4F5B", x"4C484646", x"54754441",
									 -- x"41444B38", x"4E4D564B", x"3A4A5D70", x"654D3C45", x"3D353740", x"4C2D3233", x"36213D49", x"38423A42",
									 -- x"3F363940", x"3E3F423F", x"3E3C4244", x"3D2E404B", x"3B425348", x"443A4247", x"44573D2A", x"3A38423F",
									 -- x"382C3B43", x"555D4943", x"63404661", x"4F4C645A", x"37313438", x"35353B2A", x"38433F3A", x"383A303E",
									 -- x"3440413C", x"2F374D56", x"4A3D4836", x"43273843", x"3736331F", x"435B4D48", x"3C263E43", x"393E3832",
									 -- x"3B35343D", x"41383846", x"443A4741", x"3A4A4938", x"2D42402C", x"2B474936", x"47494E47", x"434F4A3C",
									 -- x"3B283948", x"3F483F38", x"4D4B443A", x"4835303B", x"2F3A4849", x"463D4D42", x"47443E36", x"443D394A",
									 -- x"503D5144", x"453C4E46", x"5F444548", x"36363640", x"37433B40", x"4430343D", x"38424A46", x"3B494149",
									 -- x"44404449", x"4A56434C", x"3C4A4C58", x"584C4B43", x"3B3B3544", x"54413F4A", x"43555760", x"695A4655",
									 -- x"65585952", x"7357415A", x"515F6460", x"55625655", x"524E604B", x"4B4C5755", x"50614C5A", x"584F5960",
									 -- x"4D50634E", x"47674D4B", x"5C526056", x"534A5B53", x"53594C54", x"4C566036", x"48425248", x"423A4035",
									 -- x"3C4D4B4E", x"45454B5C", x"685C535D", x"544D3853", x"3C4E4D42", x"44474E38", x"4B5F4C4F", x"543D4841",
									 -- x"3E485D53", x"565A6164", x"44495F5A", x"5B425161", x"696A6996", x"8D977C62", x"6F946378", x"7D61707E",
									 -- x"7D879295", x"96777B62", x"71696148", x"5C50724B", x"53465C61", x"6649505B", x"455C5843", x"575F4454",
									 -- x"4F413953", x"4F4D3955", x"454F5A4A", x"453A4E50", x"52707A83", x"726D7264", x"60686254", x"6E6E5E6C",
									 -- x"756A6954", x"514B5F6C", x"65937A6A", x"78668168", x"69737E74", x"6D757978", x"79647675", x"73637677",
									 -- x"746A6F65", x"655F5A75", x"5A585A68", x"64665358", x"65524F4E", x"715C5E63", x"6B746B61", x"56586E6F",
									 -- x"50534A42", x"4646464F", x"53504F49", x"56725645", x"575D5946", x"4A515047", x"4F434146", x"37434D36",
									 -- x"755C3E54", x"66676B44", x"575D616B", x"7C566083", x"5D66525D", x"79686659", x"6B726D78", x"6B7B746A",
									 -- x"6B596365", x"565B5A64", x"60595254", x"625B4055", x"6450494E", x"5A484749", x"4141494E", x"46424857",
									 -- x"5A534F41", x"4C4F5847", x"574B483A", x"3D444347", x"3C55634C", x"51353E53", x"47484047", x"432E4F5A",
									 -- x"4A4A5052", x"4C544147", x"3F494C3E", x"51403B3E", x"3A304838", x"221D3134", x"34393640", x"383B3936",
									 -- x"3D332F2E", x"292B3D51", x"443B5C56", x"48373949", x"46673435", x"413B3C42", x"41424E3F", x"414A4259",
									 -- x"2A383E38", x"3D313A31", x"2B162B36", x"3753484F", x"39353E3E", x"3125393D", x"3E474E42", x"3B30383C",
									 -- x"46352437", x"414A4E51", x"5449453B", x"3A293343", x"284B3632", x"48514131", x"443A384E", x"4435333A",
									 -- x"31393932", x"36434642", x"47344147", x"38363B40", x"47443B40", x"3F433D3F", x"4F454947", x"433F3F37",
									 -- x"39472B43", x"40444844", x"4C505040", x"4A4C4B3C", x"49423C42", x"4A41434A", x"49233250", x"503E3C35",
									 -- x"37453C38", x"4F4D425C", x"52425358", x"545A4C44", x"3F3A3B42", x"412E3939", x"2A45413C", x"413A3733",
									 -- x"25405044", x"27433648", x"3E494951", x"51413D44", x"43494137", x"373B4835", x"4B5B4337", x"42423E4F",
									 -- x"4F5C4A53", x"4D514439", x"393B4844", x"445A3F66", x"44354250", x"53504641", x"3E53434B", x"344E523F",
									 -- x"3835444C", x"4C525645", x"42436052", x"45576667", x"504D5355", x"485B624D", x"37574E4E", x"4D365133",
									 -- x"5B634F51", x"4F535457", x"54525350", x"4A75524D", x"4D6D5359", x"59526855", x"584F5D6E", x"604F595F",
									 -- x"616B7D62", x"5C476267", x"7162615F", x"755D595B", x"625D6394", x"7F7B7F68", x"78977C73", x"9271706F",
									 -- x"7C645353", x"555E6A49", x"54565E57", x"6F515658", x"4B54492F", x"382C484C", x"58603D39", x"42455952",
									 -- x"3E38324D", x"3F343645", x"48544C3D", x"5058554C", x"5964705B", x"5B5C4C4E", x"4D354737", x"4D4D5A5D",
									 -- x"615D6755", x"5C564F58", x"68355466", x"66656968", x"7A816D65", x"6E75697C", x"825F6B7B", x"8273655F",
									 -- x"736E686A", x"5E615C66", x"6C636366", x"6475BF76", x"63DFE2B7", x"5F6E6D5F", x"68837B72", x"67585F62",
									 -- x"4E454D51", x"46484E45", x"504C4E51", x"4F523F49", x"5A4F4A4C", x"465B4A58", x"4B474844", x"4144534A",
									 -- x"583D495E", x"5F5C5F61", x"6E697783", x"6B59667B", x"78637575", x"70625F61", x"68657969", x"5F6F535D",
									 -- x"55415E52", x"464D4449", x"5E506270", x"585C5F5A", x"4C404B48", x"302E4531", x"3F324B4E", x"56553943",
									 -- x"6356504F", x"444E3A40", x"52475449", x"3E474D45", x"4E455651", x"514B4C4C", x"5A554E57", x"4A5C453F",
									 -- x"45663E5C", x"44343241", x"523D3A32", x"40393D31", x"27363C41", x"433B3C3E", x"311F4545", x"1F2A3039",
									 -- x"182F352E", x"2F32343B", x"3B343F2D", x"2A35343A", x"4F3F1534", x"3E4D593B", x"3B514840", x"42523B31",
									 -- x"3442313A", x"373A3A36", x"38453F4F", x"3F454042", x"2A44473F", x"4B3F3938", x"353A4747", x"3C354B44",
									 -- x"40474146", x"4144474A", x"4D5B4A48", x"40484D4B", x"4F663F35", x"3B3B3C3B", x"303B3C45", x"38393936",
									 -- x"3D363334", x"3535393C", x"2E3A3E2E", x"2D43473A", x"4444414A", x"474A4C5A", x"463F4645", x"49404741",
									 -- x"4550554B", x"453C3F4E", x"55505744", x"324D664F", x"60474452", x"493C3E51", x"453E3F42", x"37424C45",
									 -- x"393B413A", x"294F5B4A", x"523B3833", x"44554741", x"36372C2D", x"49392B38", x"253D2B2F", x"3C1F543A",
									 -- x"3740274F", x"3A3E404A", x"4146443F", x"4B4E4043", x"43433746", x"2B303742", x"2C523C39", x"324C4048",
									 -- x"50604F49", x"443E314C", x"39373B3F", x"452D413F", x"47565A47", x"3C464337", x"51434A6A", x"59534A57",
									 -- x"68525771", x"53506459", x"596B595D", x"5F6A5B63", x"5C638361", x"7F706F6C", x"567D7561", x"605E6B6D",
									 -- x"57625356", x"595E5A4F", x"56454354", x"4D513B68", x"55615D4B", x"4A624D57", x"5F525C5E", x"545A5C5E",
									 -- x"53606277", x"5E555D57", x"8B645C61", x"6A6B776E", x"59666666", x"70495961", x"666B657B", x"6B656265",
									 -- x"7D6D5C61", x"63685C57", x"5965535A", x"554C5A73", x"5F616451", x"5D4A2C36", x"4D521B29", x"0E1E4242",
									 -- x"494D4F3F", x"51554942", x"4B5A6461", x"65666F7B", x"4F5F6F4A", x"4E453049", x"5B384D4A", x"555D6D69",
									 -- x"60526363", x"535C3B3B", x"4F514256", x"5D596A52", x"67687066", x"55495E79", x"645E555F", x"5C69664D",
									 -- x"615B7166", x"5E7C706B", x"7F696174", x"7251D5B2", x"44FFFFFE", x"3D347A71", x"6B6C7A8B", x"7B5F5B60",
									 -- x"494C575A", x"504B4C4B", x"4B4C5257", x"4D3C3D5C", x"47283C4C", x"43595B68", x"55455A64", x"55537065",
									 -- x"64776370", x"615E6B6E", x"6B706673", x"5A766152", x"6C72686A", x"5D5F5463", x"6D4D3E5A", x"58605655",
									 -- x"57545645", x"47454A4E", x"54665A45", x"59595448", x"384C4F5C", x"46434E59", x"585A565C", x"60575078",
									 -- x"6058584B", x"4D5F4B54", x"434E524B", x"53524A4C", x"3748544F", x"3A43444B", x"45495A48", x"34373618",
									 -- x"313C402E", x"332E3E31", x"3B3D3A3A", x"373A3634", x"23393C53", x"3E345B50", x"4F4C403B", x"27192E32",
									 -- x"1628261E", x"282D2C33", x"2E323036", x"37383E3D", x"4D463E3C", x"563C2731", x"38541F4D", x"5D40362C",
									 -- x"563B262F", x"4B564643", x"44353D44", x"29352B39", x"34423B32", x"3B3C3B36", x"3637374A", x"3839493D",
									 -- x"41453C40", x"45474139", x"3549444D", x"4B49453A", x"3E3E3432", x"35313136", x"2627413C", x"253C3A32",
									 -- x"41474438", x"36464A3B", x"403F3C3C", x"3E3A383E", x"414E4835", x"2F414338", x"333F4440", x"494A4E42",
									 -- x"4C404B4F", x"484B4B4F", x"384A5454", x"5E625E59", x"4F4C4642", x"3D413340", x"4947485A", x"46444950",
									 -- x"583D3D42", x"433D3C3D", x"4F403B37", x"443E2E31", x"453C3938", x"3B37393C", x"33373A46", x"35445B37",
									 -- x"414D2C38", x"3259553C", x"373B4241", x"4C4E3B3F", x"3743434B", x"474A3D3E", x"3E3D3439", x"3B494B54",
									 -- x"5B57483E", x"603A404A", x"43444A43", x"4C434749", x"5B5D523C", x"41435060", x"444A5759", x"5C544656",
									 -- x"60554257", x"464A3846", x"4C543C4C", x"654F6766", x"4F715E6E", x"6E68816B", x"5B796C5D", x"666A5F6B",
									 -- x"55616662", x"5D5C6058", x"4F7DB652", x"60736077", x"5C684D48", x"47B3F689", x"4B626058", x"52515460",
									 -- x"6F60625B", x"624E6C5A", x"56645F62", x"756C6172", x"5F756762", x"765E4E58", x"4B595F53", x"555E7659",
									 -- x"5A5B6064", x"57635953", x"4D506D57", x"49444138", x"5E395158", x"40556C5B", x"4D4C333A", x"32404854",
									 -- x"5D57465E", x"5D5C4F48", x"4D4B6869", x"59565D54", x"3D4F5147", x"5D505061", x"5C515758", x"53565056",
									 -- x"4E3E6B63", x"5D78785F", x"5D766A5A", x"68757583", x"5C3E6A52", x"5E585461", x"61636365", x"67548777",
									 -- x"62627A72", x"6B6A8386", x"68657F73", x"64684F68", x"6C5B7489", x"69636A79", x"644D6578", x"615D685F",
									 -- x"50534A4A", x"5753484D", x"51635D54", x"5D5D5D55", x"5C52635F", x"637F8A6E", x"747F7C75", x"6C5C5A5D",
									 -- x"5D664665", x"60576660", x"605D5762", x"6F6D625C", x"69644B63", x"3F49555F", x"51455360", x"536A5954",
									 -- x"464D4342", x"403D4C4A", x"4F6F4141", x"4D5F5554", x"446A5857", x"4B3F3645", x"4847304E", x"6B545253",
									 -- x"4348482D", x"3B453026", x"4C4E475B", x"2E393535", x"39504136", x"33405553", x"0F3E3A3F", x"3A332A41",
									 -- x"423E2E37", x"50393530", x"1C423F2F", x"283B3026", x"2A2C3E3C", x"3E3B373A", x"382F3E38", x"27213931",
									 -- x"1E201E20", x"27272428", x"2C212636", x"31273845", x"41444343", x"453B142E", x"3141485D", x"46413A2F",
									 -- x"372D3135", x"5040302B", x"443A3443", x"312A3832", x"32323338", x"2C293132", x"373C2F41", x"362D372F",
									 -- x"3A36303C", x"4C433B36", x"3B4A4835", x"31332E22", x"3238363F", x"31383E32", x"2F3A4234", x"32362537",
									 -- x"3B313137", x"383B403F", x"2E363735", x"373B3C38", x"3D383935", x"34383C35", x"33393042", x"463D343B",
									 -- x"4340344C", x"4E534E39", x"3C3E4346", x"5A473B3C", x"46565147", x"4F674845", x"5047404D", x"3D4B5446",
									 -- x"414B565D", x"444B4750", x"4F443F3C", x"41343742", x"54624D44", x"4035363D", x"3624403A", x"343C321E",
									 -- x"36353D35", x"2C413A3A", x"30383C3B", x"3D382F31", x"4E384348", x"534A4244", x"6A384246", x"50445053",
									 -- x"4A5C524D", x"4F575F3F", x"485F3E40", x"403D4346", x"3C696750", x"4B464354", x"4E4E4D5A", x"5244344B",
									 -- x"3A403632", x"54444755", x"49363E48", x"4449535F", x"54454E52", x"3E405C47", x"5163505C", x"6B5C4F51",
									 -- x"60617365", x"564B5556", x"4E76CE5B", x"394D514E", x"514B4F6E", x"6576BAA8", x"4B526054", x"58634355",
									 -- x"5D5A5D52", x"5A606458", x"5B56504E", x"54585854", x"5055585C", x"575A4C56", x"57514752", x"545E5F5C",
									 -- x"50495B67", x"544C5247", x"492D5657", x"494E3D4F", x"574F444A", x"5850474A", x"58456465", x"51565B5A",
									 -- x"63645D66", x"5E4C5E5C", x"5E63716B", x"726A5F5D", x"70644A52", x"695A645B", x"565B5955", x"58585C69",
									 -- x"59667761", x"74726C62", x"655B6462", x"5B657159", x"5778555D", x"8C585F57", x"5D5C6C85", x"67485854",
									 -- x"4B545160", x"6847615B", x"5B4A3B4E", x"545A5A56", x"59524656", x"655A605F", x"61696A66", x"6768635B",
									 -- x"534E5053", x"51525859", x"606D6C73", x"785B5D63", x"6B736D7C", x"66616365", x"39616259", x"5458575E",
									 -- x"5C4B6561", x"59675A45", x"54585265", x"5863706C", x"5C3E4949", x"435C604B", x"58655F61", x"665A444D",
									 -- x"4D494D58", x"40434E42", x"48684B49", x"482F3F56", x"53524B54", x"452F3839", x"46414C3D", x"493D4D40",
									 -- x"41493230", x"3B4F3B40", x"603C2B38", x"33323924", x"413E3A3D", x"3E30644B", x"41474A4B", x"44322433",
									 -- x"49182D41", x"24243C53", x"4F322B32", x"323C4D50", x"3F2D3638", x"341F323B", x"30292325", x"271A4950",
									 -- x"36343028", x"25303832", x"28123037", x"312E2E32", x"413F3D26", x"36333540", x"363D3A3C", x"36363237",
									 -- x"3445313B", x"3B2F2C28", x"2F394442", x"3B2A3029", x"2A332423", x"1E1D253D", x"2B362C33", x"3A212F2F",
									 -- x"39352A24", x"2E283541", x"3C3C4234", x"323C3B49", x"2D4A3242", x"1A364E2E", x"2A333534", x"2D2D3533",
									 -- x"3026272D", x"2D313633", x"2F322F29", x"2933311A", x"33313F3F", x"3A353E39", x"384B3442", x"3D422F30",
									 -- x"2E403A2A", x"3F3A4238", x"3C41433D", x"5F3C3548", x"5C474748", x"38564C48", x"55403249", x"4D4D4E48",
									 -- x"4A4E594A", x"55504C43", x"483B3739", x"423A3F3C", x"43533D46", x"40373826", x"4E403A50", x"5A3A4B69",
									 -- x"45364453", x"5E4D4537", x"3A493B2E", x"37495345", x"45314544", x"2C434137", x"52284048", x"3F444F4B",
									 -- x"4B415D4B", x"47584F48", x"4A463E3A", x"34394848", x"43654A4D", x"5052364C", x"514B4170", x"5152424C",
									 -- x"47453B55", x"614D5C3A", x"5F564A4E", x"4F4B4337", x"45234A50", x"3B453E4C", x"50524C59", x"5F4B4657",
									 -- x"584D6961", x"574B575B", x"61533957", x"4653525D", x"7251504F", x"604C3D36", x"585D565D", x"6571604A",
									 -- x"5C5F6446", x"5A6B5648", x"4948585B", x"5A5C5D47", x"533F6159", x"6556555B", x"6F46575D", x"555A5552",
									 -- x"40525751", x"5341524B", x"68565652", x"504A5063", x"6A575B41", x"4A4F3A4B", x"4A495765", x"616F5E70",
									 -- x"656D7970", x"93907383", x"8D656E71", x"72686C68", x"6D6D7685", x"785A6F6F", x"67656D63", x"77697267",
									 -- x"6C664F69", x"5B5A596C", x"675F6560", x"65535451", x"66626A68", x"5C4A3843", x"65576B63", x"4152463F",
									 -- x"3F53494D", x"5C56524D", x"56605954", x"564F535E", x"5F5E5262", x"4F3F5367", x"5F625F5F", x"595C6352",
									 -- x"66626967", x"5D676E5B", x"626D635D", x"7659675C", x"5D606058", x"414A4C41", x"4C4A5154", x"555A6A5E",
									 -- x"5D4D5951", x"5C65585D", x"594A545A", x"54635C3C", x"5467514D", x"506A4F47", x"5450594F", x"4A4A454D",
									 -- x"5A4C5665", x"37454141", x"45644457", x"52566261", x"5F4A496E", x"4E5B5C4E", x"6B60392A", x"3F414149",
									 -- x"4748454E", x"187E663C", x"4324373F", x"43353322", x"3C483932", x"34493F2A", x"3433404E", x"41434244",
									 -- x"3C3E3D44", x"4A474745", x"45374649", x"413C4235", x"31303530", x"2E294247", x"352C2E28", x"28404633",
									 -- x"2A3B3C3B", x"324D3A4B", x"343B3A35", x"31333133", x"35373A32", x"2E2D3A3F", x"553A3039", x"28303637",
									 -- x"443B232D", x"26302A2B", x"253D333E", x"3519092F", x"2F242E30", x"212D3B51", x"31241A23", x"2126302C",
									 -- x"461A3E2A", x"2F373B49", x"343D3337", x"3131363F", x"4241453E", x"442F4634", x"3126332A", x"35353426",
									 -- x"1E293D42", x"323D3933", x"30352F24", x"3C37312E", x"2F2C2E3A", x"3F313D33", x"30403C40", x"40323641",
									 -- x"3C4E4F46", x"4C3E3E40", x"3542463A", x"45383342", x"5A3E3030", x"39443643", x"3F3F394A", x"4A4F4E3E",
									 -- x"42332D4D", x"4F414429", x"31314348", x"3A352237", x"40363F4A", x"3C4C3540", x"3A3E3039", x"484C4352",
									 -- x"4239412E", x"38404843", x"45495343", x"4449324B", x"45455B48", x"524F5947", x"45474D43", x"4B566B4C",
									 -- x"4B65474F", x"3E464243", x"3B315747", x"3A535F51", x"4038384C", x"55626A58", x"413A5F69", x"534B5A63",
									 -- x"695B556A", x"585C796F", x"54664D5E", x"7A4A4140", x"493C5C73", x"5759585D", x"50654849", x"545D4D55",
									 -- x"4F555249", x"40384E54", x"5C674D4A", x"565C5C52", x"4F315361", x"594F505D", x"5B5B5E5C", x"5B5F6C56",
									 -- x"2C4C623A", x"44435354", x"5E4C5059", x"56595B57", x"655C5349", x"655F5D77", x"5A52787A", x"5B545C52",
									 -- x"574A534C", x"4745512E", x"4C555363", x"3B4E4D4D", x"6050475E", x"65616658", x"545C5958", x"5B6A6569",
									 -- x"59696370", x"72737774", x"79545C5C", x"646E7173", x"597F8E81", x"7D7E6E6C", x"82746A91", x"77797F77",
									 -- x"6E777A6D", x"757D6C97", x"7365837E", x"8A7F7888", x"8276766E", x"7246645F", x"656E5658", x"4E4A5832",
									 -- x"2E5B4F3D", x"4242505F", x"6E7C7A82", x"62615C65", x"8C675F59", x"645D5B70", x"6B586467", x"4A5B615B",
									 -- x"5F656A6F", x"6D606275", x"6C5E3A4A", x"6B5C5B45", x"4C4F5651", x"50404A5C", x"646D6659", x"596F5861",
									 -- x"5D5B675B", x"5352484E", x"474A4B55", x"5D70674C", x"4F53544F", x"4A363E3D", x"394C5845", x"4C485347",
									 -- x"47244E4E", x"543E4644", x"3936444A", x"50664055", x"5551442D", x"3A38515A", x"34332136", x"60403D41",
									 -- x"36543C25", x"3754472F", x"3E5D4140", x"443F312D", x"3F432E4E", x"D2FF9A11", x"403D474A", x"46464A4B",
									 -- x"36384643", x"3C515330", x"304B5140", x"4B3D2E3F", x"393B4D3A", x"4A404A3F", x"2727413D", x"393C3827",
									 -- x"30393642", x"383C3242", x"45453A3F", x"34473331", x"2E2F2E3D", x"2B34333B", x"39353B33", x"383C2350",
									 -- x"42312F2C", x"2B2B4229", x"25342F43", x"2E252A39", x"34302E43", x"4A49313C", x"290F3253", x"282F2832",
									 -- x"3A2E2C41", x"3337413B", x"363B3137", x"304D3949", x"45343E33", x"313E373B", x"32305440", x"413C363B",
									 -- x"35374F43", x"3D3E3B38", x"1617303F", x"46253239", x"31372D44", x"40403A2E", x"312F3637", x"4047303C",
									 -- x"3D474340", x"3E403F37", x"3F463D42", x"483A3841", x"3F433A35", x"34463B44", x"4048513B", x"333D3644",
									 -- x"3E273945", x"3A384037", x"383A4245", x"3E3F4C35", x"40442C3B", x"3236333C", x"49334A59", x"2A38492B",
									 -- x"3C304539", x"2C4C474E", x"4E4E4645", x"4A4B5B46", x"3941394A", x"5B324252", x"423A4A46", x"42524B3C",
									 -- x"4D4B3C51", x"464B3E3B", x"3F3D4B43", x"48515551", x"575B574F", x"57606367", x"545A7540", x"4E595756",
									 -- x"5D536957", x"4C596155", x"434C4745", x"3C425C5D", x"4F5D5B5C", x"5F605B61", x"6D4E5561", x"52555354",
									 -- x"60674F50", x"4F525B68", x"40563B46", x"59324D48", x"4B3E535A", x"55556568", x"47625047", x"52504E69",
									 -- x"34454036", x"40314F56", x"5B624850", x"5E5A5749", x"55585359", x"68654C57", x"58415A5F", x"5C55463E",
									 -- x"54515150", x"4C544A41", x"48456F43", x"4B7E5866", x"5A5F7250", x"5A565678", x"7E5B4C4C", x"614D5659",
									 -- x"6068575F", x"584A5C4D", x"5A716066", x"76705C84", x"64666F7C", x"7E7B6E72", x"9F705873", x"60657A70",
									 -- x"6E6B656F", x"6C6D5263", x"67736570", x"7F969B7C", x"8E9C919D", x"95736A7A", x"887F6A5B", x"615D8082",
									 -- x"6973716B", x"78635D5B", x"6468545E", x"656E6E70", x"6D817863", x"77867482", x"81847675", x"585F6662",
									 -- x"58607076", x"695C5F69", x"595F565E", x"59565862", x"58506A7A", x"725C605F", x"544B5954", x"6A594652",
									 -- x"564C5D47", x"42504556", x"535A5142", x"6974744B", x"59797853", x"51504562", x"5E58616B", x"454A4234",
									 -- x"2F405540", x"5149343B", x"39453D30", x"3E264952", x"69865438", x"3E624C3F", x"3B47494B", x"2C463B3F",
									 -- x"442D3C49", x"254A413C", x"43533F36", x"4F424847", x"3F433846", x"79922628", x"45495249", x"453C4952",
									 -- x"3E464F48", x"484B4040", x"52614253", x"4A2D3647", x"4F343841", x"333E3A44", x"4D494B4A", x"30413135",
									 -- x"232A2936", x"2F2A2D37", x"21243621", x"2431322F", x"2B2C321B", x"30283736", x"2E323C3D", x"37223252",
									 -- x"432D2741", x"2B243E4A", x"48465437", x"2C5B5229", x"37393661", x"4B31292C", x"34204527", x"53453A2B",
									 -- x"3C2E2E3D", x"3933331F", x"26383F37", x"35413541", x"2C312D30", x"2E3A4037", x"38384E39", x"3E303137",
									 -- x"3C383738", x"302B4532", x"2B3A372A", x"2B3A2F43", x"36483837", x"2E3B3A31", x"373E373B", x"3D3C3639",
									 -- x"3F464348", x"424F4D3C", x"393B2842", x"433C3B3E", x"31424041", x"4E5B4D45", x"48403D42", x"3D2B2A31",
									 -- x"3F3F4437", x"3B3E474F", x"3E243E34", x"3A3A4142", x"49534B57", x"53543B49", x"4237393D", x"42403E33",
									 -- x"40365356", x"52434F38", x"474E4941", x"4B3F6845", x"45411332", x"453E3E40", x"3E423B42", x"34425C5E",
									 -- x"3E407044", x"47484B4B", x"4F4C2E40", x"433F2B49", x"5F435850", x"52544B50", x"573F5E54", x"3F2D5B5A",
									 -- x"4B67704B", x"44535C55", x"59625B58", x"48696560", x"6F605B5F", x"6E56445B", x"4F485051", x"514D5357",
									 -- x"4A28464D", x"60504A5B", x"58544C59", x"59535E43", x"454B5351", x"4B4C533D", x"4732413F", x"514F2849",
									 -- x"4952483A", x"474B5253", x"5647374D", x"5F553B42", x"3E585A4E", x"6C5F4C5C", x"595F4B58", x"575F5F51",
									 -- x"5A405670", x"58524D54", x"415F6048", x"547D4C5C", x"57557E44", x"544C4B5C", x"68523C47", x"574F5255",
									 -- x"60675635", x"575E515E", x"5F695861", x"84765F62", x"666B5677", x"78835968", x"6D6F4A85", x"8D5C7463",
									 -- x"5D66566F", x"6F716F5D", x"53747270", x"6F708556", x"6A737877", x"7A756681", x"B29E6D73", x"84556974",
									 -- x"70747073", x"72736C66", x"6F8F6752", x"546E666C", x"686D8771", x"8872706F", x"819F9C77", x"7C686871",
									 -- x"5755564E", x"42465151", x"5D5A6261", x"60755D5E", x"645C6771", x"5658594C", x"3A504E4B", x"413E424D",
									 -- x"3939493F", x"464B4C4F", x"564B3153", x"5D574E4E", x"5869544F", x"42556864", x"54496346", x"2D4E5156",
									 -- x"52766A64", x"58664553", x"4E504247", x"5F6B5E51", x"4B40433E", x"52344657", x"45314762", x"44423A4E",
									 -- x"43574955", x"6C4C3F54", x"49324F6C", x"4B43586E", x"4A3D3A45", x"3242505E", x"4C4A494B", x"504A5258",
									 -- x"4D385567", x"5D564947", x"45464C3F", x"40403B39", x"31173B36", x"2138362B", x"4D49403B", x"20392B3B",
									 -- x"343C3D33", x"25242927", x"2B33402D", x"203B3131", x"3E373336", x"67504146", x"455A4B41", x"39595043",
									 -- x"555E4A52", x"46615248", x"454A5248", x"44496748", x"583C3164", x"3A321F39", x"4D31321C", x"38323B2E",
									 -- x"43343931", x"2D273632", x"3D4B372D", x"35323C39", x"2E2A3324", x"2F3D3428", x"39392F30", x"46313928",
									 -- x"322E2E34", x"34423C3E", x"2E3A3B11", x"2F413139", x"34221A2B", x"432F2F32", x"303E393C", x"3E343E3E",
									 -- x"434B484C", x"494D4636", x"41402E4A", x"3F403737", x"2F3C3C35", x"3E35373C", x"2B453B39", x"3631373A",
									 -- x"25495041", x"3F333D34", x"2F3A3A24", x"2E233434", x"3B424451", x"4F5C4658", x"45353526", x"424F532D",
									 -- x"42342747", x"443B4B41", x"655D3A33", x"37444A45", x"4E44413C", x"46405A32", x"3E463C49", x"5050664D",
									 -- x"44444A35", x"464B3F43", x"4B565234", x"53424459", x"4F5F5463", x"3C3B5753", x"4E513143", x"66585552",
									 -- x"5B794F58", x"6061675A", x"51576558", x"6164645A", x"3F3A6064", x"615B5C54", x"626D3933", x"564D4E4C",
									 -- x"574F2342", x"635A4D47", x"39354C4E", x"4A5A5A42", x"4B484647", x"484B4C3C", x"4A4A4248", x"3C4B4738",
									 -- x"4A64424E", x"6F6B6E78", x"75517247", x"3D6F3E55", x"4750474B", x"384C4548", x"4E4B514E", x"51725F5C",
									 -- x"4656615E", x"635F6B86", x"7967557D", x"5868443F", x"4A504E43", x"4757535A", x"4D655454", x"5D625265",
									 -- x"513C543F", x"6273595B", x"665F6764", x"6D6C7466", x"66777A51", x"445A5D41", x"6E6D577A", x"90747184",
									 -- x"6472576D", x"726E9187", x"7D767668", x"635F7060", x"6A756563", x"5A556759", x"5D404E69", x"5F5F6C6B",
									 -- x"54747465", x"645B6C7B", x"8D7E7E7F", x"68666A7A", x"696E6B6F", x"526D6564", x"7687A978", x"7355536D",
									 -- x"535B534F", x"5752484E", x"575A605E", x"5F695A55", x"5264645B", x"4B4D4543", x"50655448", x"45423D44",
									 -- x"4B51453A", x"402E4D44", x"514D5573", x"6D52616B", x"69434F5E", x"5C5B5255", x"3F3F3F2E", x"54734F58",
									 -- x"70545266", x"53464E4F", x"4F6C4954", x"5E444E2C", x"473F2E3C", x"3C463B2E", x"3F60434C", x"484B5350",
									 -- x"586E4B6B", x"3B473F42", x"3F1F4468", x"4A485E62", x"515D5659", x"375D5645", x"4D3D2B40", x"504E4540",
									 -- x"2F355244", x"252A3544", x"3A2E6551", x"433C6234", x"2F224A56", x"364A3544", x"433E4124", x"262C3038",
									 -- x"303A4A3A", x"3544484A", x"4037413C", x"40524141", x"423D3E44", x"5C483F46", x"50794E48", x"70555057",
									 -- x"6D596461", x"5F4E536A", x"56505456", x"49303647", x"484A7533", x"44443B3A", x"2C352F35", x"32362B38",
									 -- x"332F232F", x"2A25382D", x"3347313D", x"3533302E", x"30272426", x"3630200D", x"33372B3B", x"533F4331",
									 -- x"4053313A", x"3F2F2F34", x"37322439", x"29202134", x"36343624", x"2E1E323D", x"342C3C30", x"3C393233",
									 -- x"35474A43", x"43363A41", x"44464051", x"414D3F40", x"3F463E3F", x"3C34333D", x"45523F29", x"354E3B4A",
									 -- x"3D393E3B", x"2E324123", x"2F3C3D35", x"433F484D", x"43493747", x"363A3B3D", x"2E373E42", x"5F513C30",
									 -- x"634B3237", x"4047485D", x"57444A46", x"62545653", x"4F3E3062", x"44405D49", x"46404F39", x"4D525A44",
									 -- x"627F4D4A", x"5F56514C", x"574F6651", x"6B484F7B", x"4D5E5469", x"54593F55", x"3D484C55", x"5E685C5C",
									 -- x"635D496D", x"68616055", x"4E535B61", x"56535846", x"5D403F4C", x"4B4B754F", x"514F2B3F", x"4625314D",
									 -- x"4B664F4B", x"2E3F5850", x"4B532F51", x"435B3545", x"5D535357", x"58544949", x"4B543D51", x"3E493F59",
									 -- x"6B394F65", x"494F4D5D", x"5A545E5C", x"596C5E53", x"484E4B3D", x"454B5859", x"4E484C4E", x"38474B4F",
									 -- x"485A5865", x"77545467", x"62525F4E", x"394C2A38", x"435E4A4E", x"5C595767", x"6B5B767B", x"6069766D",
									 -- x"71566971", x"775E535A", x"65626055", x"48636264", x"63758172", x"80756D6F", x"6F6E736D", x"585C5462",
									 -- x"6B4D606C", x"787F5376", x"81767270", x"5857484C", x"61545D51", x"40665C67", x"64543F5C", x"604D626F",
									 -- x"75936767", x"736A6780", x"726A8A79", x"756A616D", x"6A535E58", x"70607077", x"77667E7B", x"686E6E75",
									 -- x"5256534B", x"494D4E4B", x"50564854", x"594C5450", x"58595748", x"49495150", x"4A25494D", x"4547482E",
									 -- x"403C4B44", x"56505652", x"4B646375", x"4C626764", x"5A594A5D", x"51474850", x"5B635057", x"5C5C4459",
									 -- x"54384348", x"483A5652", x"504B432B", x"4E2B4030", x"494D4750", x"4E473F40", x"39645264", x"5A6A635A",
									 -- x"565D3D39", x"5E5E5B68", x"485E5D4E", x"4D4F7579", x"44326D48", x"3F4B4539", x"3636304B", x"4D4C5156",
									 -- x"42545B4E", x"53554341", x"45483E53", x"69565C2E", x"3B406323", x"31393A3F", x"4D453A23", x"363A3C3A",
									 -- x"2E334538", x"37423A40", x"44384C44", x"513E3B4B", x"5642484A", x"3C334C5C", x"4C446949", x"43424A54",
									 -- x"7151624C", x"45394A43", x"53444B43", x"3F57243A", x"5F4C4A3A", x"43394448", x"2F344539", x"35332932",
									 -- x"3E313837", x"3B2D2F25", x"2730312D", x"23262C38", x"302E1129", x"30223132", x"37323132", x"332F323E",
									 -- x"2E223737", x"322E3437", x"2A124244", x"4E3C2A50", x"2F2C323D", x"42363B48", x"3D31332C", x"352E302E",
									 -- x"3E3A2925", x"3F3A3835", x"32373B40", x"36473F40", x"3B3E2F3B", x"2F3F3239", x"403C3C40", x"3945494D",
									 -- x"31172733", x"333E342E", x"573C4D4B", x"4B503941", x"3C393A45", x"313F353C", x"1F192F4F", x"373A3524",
									 -- x"49504038", x"4D3E3F50", x"47473C6B", x"474E434C", x"564F6D5F", x"324C4858", x"69646D49", x"5558726E",
									 -- x"375A4C3F", x"56585A62", x"55484C46", x"4A50435E", x"4C4F5649", x"5F4D5A65", x"70514A64", x"806C6056",
									 -- x"5F436B6B", x"4D646256", x"5C675458", x"4F4B4E42", x"6C4D5B47", x"5D7E7251", x"4D5B594D", x"4A57544F",
									 -- x"49414B42", x"4B503F50", x"4446604A", x"52332B43", x"3C4D554E", x"4E584C47", x"3947684C", x"5062526F",
									 -- x"4C4C565F", x"46484951", x"43515E50", x"50585255", x"5A41507E", x"5440608F", x"55574F43", x"4235704D",
									 -- x"40606362", x"49364A48", x"494B5141", x"393C5956", x"39443B4B", x"50524847", x"4C4D5057", x"56615755",
									 -- x"59586660", x"5642395C", x"5B596A5A", x"4B616364", x"686F7285", x"708A7971", x"647D836E", x"58717167",
									 -- x"6E8D5774", x"5F384A58", x"6B6A5F68", x"787D5C43", x"6C617061", x"6275626B", x"8F646567", x"7C7F91A9",
									 -- x"81706A7A", x"7278845E", x"6C626766", x"68815E5E", x"75666F78", x"8987887E", x"788A867E", x"8189927C",
									 -- x"4B49595B", x"494B5244", x"4751444E", x"50414851", x"5B535B5C", x"5E575547", x"34424743", x"435B4D5C",
									 -- x"5546534F", x"595E5053", x"58555351", x"3F475251", x"524C4641", x"2449535B", x"54505F56", x"51434F3B",
									 -- x"313F4B3C", x"45534F56", x"4D4E584F", x"6058494A", x"5354544E", x"554A5456", x"50475D57", x"5E616458",
									 -- x"624C3448", x"7C557B4A", x"5A784442", x"3B5F595A", x"315C6343", x"3A343643", x"3A44474F", x"3E33454A",
									 -- x"3F2F3749", x"48404042", x"3C486363", x"5A6B4044", x"52405131", x"32372D42", x"3C3F2D31", x"4447413D",
									 -- x"474E514C", x"4D4F4040", x"40474A4D", x"4944405E", x"573E385C", x"4742425C", x"3F433E44", x"39453652",
									 -- x"3C44534F", x"3B405646", x"3E41364B", x"40473D39", x"2B323346", x"36103525", x"2B3A2416", x"2E28265C",
									 -- x"382A422D", x"2A19212F", x"27283329", x"2D283226", x"22223337", x"3F3D303E", x"362A2427", x"1A212438",
									 -- x"2516354C", x"3C2F3B24", x"555A3E42", x"43292D2B", x"2A353633", x"2634383D", x"32322530", x"2D253637",
									 -- x"2E352D24", x"22202930", x"2E33302B", x"2B303430", x"31313131", x"1B2B2A38", x"3E3C3941", x"453B401F",
									 -- x"2C2E3A3E", x"3A40385F", x"42434539", x"3B474233", x"3D313D34", x"253F203B", x"463C3B32", x"143F502B",
									 -- x"1E412942", x"443D3E5D", x"3C414067", x"56534744", x"514B387E", x"56494353", x"5B57504A", x"4D464A42",
									 -- x"503A3B57", x"5455444C", x"63444546", x"5B565361", x"4B48703E", x"6D657262", x"5C626E68", x"6048664F",
									 -- x"66526158", x"486A6752", x"53524634", x"503A5451", x"53655057", x"62435755", x"605A6354", x"4A464A55",
									 -- x"5231224D", x"4F4F4D42", x"3E2E4A2D", x"3C465159", x"5064574C", x"4B555450", x"545F7D59", x"4C2C4A46",
									 -- x"38475E53", x"415C504A", x"33445A6B", x"5C375873", x"5C564D4C", x"6464624C", x"646B595A", x"326E4F32",
									 -- x"4D49495E", x"6B535753", x"4A4B2647", x"62305356", x"55543855", x"30554A34", x"46563E46", x"525E5441",
									 -- x"404F6B62", x"48605963", x"5C3C4F54", x"5C6B7250", x"4A555E73", x"6A685867", x"71748671", x"75937252",
									 -- x"6B955C72", x"7659775E", x"70796C5D", x"797D6E6A", x"5E496954", x"6276543F", x"7C8A7E5A", x"63647578",
									 -- x"68769C81", x"AF8A8774", x"76685962", x"55AB965A", x"8F756177", x"77787075", x"74A0A487", x"866B7C6B",
									 -- x"574B505E", x"584A5062", x"5A56504E", x"5961454C", x"56625553", x"544C3A43", x"5E443C41", x"4343544F",
									 -- x"4A5E4F6C", x"634D5548", x"4E4F4A43", x"36484C50", x"514A3D40", x"5B4D4345", x"462E403F", x"27243546",
									 -- x"4944524B", x"49502C39", x"44525246", x"57505147", x"514D4C3B", x"424E5328", x"4446494A", x"433D5A76",
									 -- x"5E535C7A", x"4A4B7D5F", x"5D5D5065", x"586F514D", x"445D4B32", x"343D3837", x"42403E43", x"47455746",
									 -- x"48342743", x"51312949", x"4F3E6046", x"4C411449", x"572D4548", x"3E48424A", x"434C443C", x"4D3A4951",
									 -- x"4F5E5250", x"5457483D", x"54503F28", x"3F3A3432", x"35546240", x"4632302C", x"31394E33", x"414E573D",
									 -- x"4548333B", x"39314A48", x"3B3F4251", x"44425B3F", x"39464338", x"3936413E", x"39482611", x"28273725",
									 -- x"1A1E1635", x"33292D28", x"2A3D3030", x"1A193223", x"322F2E13", x"2C2C3024", x"2A231736", x"3034302D",
									 -- x"42353640", x"42412B34", x"401D282D", x"382B2F27", x"3428242D", x"2D37312C", x"2D252733", x"252B1F2B",
									 -- x"25282226", x"222F342D", x"34392D28", x"322E3F37", x"2117363B", x"3B352D2C", x"3139433D", x"663F335E",
									 -- x"38464655", x"46463E46", x"3B3D5030", x"3C4B3B59", x"3D434342", x"3A472C43", x"53513F2D", x"3E413D38",
									 -- x"3E424549", x"4C373062", x"36404E3E", x"4D393D4E", x"684B577C", x"59493947", x"674F4C47", x"38483655",
									 -- x"483B516B", x"5127583D", x"414A4748", x"48514D4E", x"46646562", x"6A3D5182", x"3B48805C", x"42698C55",
									 -- x"5B643150", x"4E474D4C", x"6E4F365D", x"59604D31", x"4F6E6E56", x"5C504957", x"4B425252", x"585C683F",
									 -- x"41475141", x"4E57745B", x"354D3E4D", x"53595447", x"4D4B3653", x"5B494C5B", x"4C656F57", x"4A515932",
									 -- x"48414359", x"52555856", x"433A3B43", x"3C33634C", x"274B5650", x"5D686A52", x"4A546E4D", x"385C5047",
									 -- x"75486466", x"5D486E5A", x"59556F5A", x"64484F42", x"253F4345", x"4D53795D", x"55614741", x"67566C52",
									 -- x"537D5E57", x"4F5E5251", x"6A545362", x"4F596456", x"645B4A62", x"4F674F4F", x"5C586772", x"66698250",
									 -- x"6D799973", x"75676874", x"6875717B", x"96A17080", x"88786773", x"73ACB374", x"7E6D7672", x"636E787E",
									 -- x"8D7A878F", x"A09F7A79", x"7988746A", x"737D7773", x"8893724D", x"76736865", x"6D5B7089", x"7F6D786A",
									 -- x"584F4449", x"3F4C5752", x"4650564B", x"4E514143", x"4C493C45", x"553D5140", x"493B4244", x"462C4D4B",
									 -- x"4147452E", x"39464A45", x"323C333C", x"4B4E534E", x"3747444C", x"3A4D2B23", x"20354646", x"3E3F4546",
									 -- x"473E4B35", x"45423646", x"443D3F4B", x"4E4F4049", x"40443A2E", x"43484238", x"49295152", x"4E4A535E",
									 -- x"543C5A58", x"49545A42", x"48573E4D", x"4E454C49", x"4A49432A", x"465B404A", x"5242354E", x"57635352",
									 -- x"48484150", x"4926483E", x"38482C49", x"3942674C", x"394A3C48", x"4E4E554D", x"425B4C49", x"4D41605E",
									 -- x"545C474E", x"514A4546", x"6945293C", x"4F442512", x"2F434130", x"443C3527", x"51391E33", x"454A3E3B",
									 -- x"3A352731", x"363B393A", x"47464344", x"3B40411D", x"2D353239", x"34383635", x"2D3E2C26", x"372E2D12",
									 -- x"492F2025", x"501F3332", x"1F262725", x"322F2532", x"40261A22", x"1B222524", x"27215548", x"2D454E2C",
									 -- x"55453A3F", x"39544428", x"162A3D08", x"312B2C33", x"352C333F", x"36473333", x"30353939", x"2E2D3035",
									 -- x"2A2F3B29", x"322E3026", x"33363A2F", x"28323B33", x"2E492734", x"2D333231", x"2C2D3D42", x"41413642",
									 -- x"53553E46", x"3B332931", x"363A3E35", x"3848394F", x"563E485C", x"435C604C", x"4B58473D", x"3B4D4E4A",
									 -- x"4445675F", x"4253465A", x"464B4B61", x"695C6741", x"575B6C38", x"453F304D", x"4B324343", x"44495754",
									 -- x"41324834", x"48583A39", x"3F525E45", x"45496B43", x"4C675767", x"634E5A4F", x"646B4556", x"57666052",
									 -- x"4B4B4F4B", x"43323759", x"66514468", x"6B5D3F52", x"594F4752", x"565B4D54", x"5B645444", x"516B5432",
									 -- x"57576759", x"5A556A4B", x"4D793B55", x"65555C52", x"3A635D4C", x"6042486B", x"524D543D", x"4B754F4A",
									 -- x"3F405A56", x"4F5A4642", x"55523140", x"536F4961", x"72605E5F", x"66795454", x"67545D4E", x"47595753",
									 -- x"514C3F4A", x"535A6B58", x"385A6858", x"7346605B", x"4529455B", x"436E7A3D", x"4843355E", x"523E4C4B",
									 -- x"5C4A5658", x"466E5559", x"5D574B54", x"515E5C6F", x"79565C62", x"49594335", x"626B6F52", x"6F8D7C68",
									 -- x"71767B8D", x"886C829A", x"766A8887", x"5F895E78", x"828F875E", x"52746851", x"5A646D5F", x"576E7B73",
									 -- x"7B72757F", x"756F7772", x"6B70705B", x"7B655F62", x"64676560", x"7D64505A", x"6973647D", x"92476D70",
									 -- x"4F4A3C3E", x"3F424152", x"49594941", x"4643494B", x"403C463C", x"44454442", x"41353956", x"4B4A4E43",
									 -- x"2B3B3F3A", x"39414D47", x"483A3E48", x"48545760", x"55686847", x"414F5E47", x"435F664D", x"484D4259",
									 -- x"424C3F45", x"3D3D473E", x"2D30444E", x"4C3A4738", x"42473144", x"42533A3C", x"43445951", x"36465252",
									 -- x"524D4252", x"58674057", x"44404841", x"4249413E", x"3E4C3F37", x"3F5A4F57", x"5432445D", x"41504644",
									 -- x"4440392F", x"2D434E29", x"404A4440", x"42442E42", x"3C3C213F", x"4741564F", x"415F5C6B", x"5B4E574C",
									 -- x"3A594667", x"484D4156", x"5B435C50", x"51433D3E", x"42484647", x"4D414B3B", x"43293036", x"3D243F42",
									 -- x"323C543A", x"3645333E", x"513E3A32", x"3F383535", x"373B3828", x"2A2E342A", x"1E323630", x"2D2F2E35",
									 -- x"421B2929", x"14223A3B", x"292F1D24", x"39353932", x"2C293148", x"2E30312D", x"2D2F3634", x"2C1E272B",
									 -- x"1C303E37", x"3A3B3247", x"3C353733", x"2F3E4330", x"48462B39", x"3A56342E", x"29313432", x"34384350",
									 -- x"302C2B37", x"32332624", x"1736303F", x"321D3D33", x"3A2E2827", x"3E372F36", x"32333D3F", x"38382C30",
									 -- x"342A332B", x"32363131", x"3E33312F", x"302B404B", x"4E3A634C", x"3E3F4849", x"34323E44", x"4650554A",
									 -- x"3B4F4D48", x"375A3F48", x"3F5C472C", x"433C494A", x"6C3A5051", x"41333D66", x"453B5533", x"404B5A2C",
									 -- x"42532F40", x"3751482F", x"26443F40", x"2F343940", x"4558342C", x"4847576E", x"5A625E4E", x"5C5A4368",
									 -- x"5355515D", x"52505749", x"212E584F", x"3560544B", x"50543952", x"3B4A3950", x"5349485E", x"4A58504E",
									 -- x"38425A44", x"453B503B", x"49655047", x"535A6D4F", x"6B53543F", x"5D463A58", x"52562E42", x"4E4C4275",
									 -- x"5F5B4A63", x"554D5265", x"5C575B52", x"6D535662", x"5853516D", x"4C434440", x"60484F66", x"4C465E3C",
									 -- x"48374E41", x"465F556C", x"633C4A66", x"5F635C3A", x"4A5F3E36", x"45535043", x"27555441", x"44344B38",
									 -- x"5B553154", x"685C5444", x"44487149", x"56446072", x"91847C83", x"6A52535B", x"6379816A", x"658D7174",
									 -- x"6C616964", x"5C595E61", x"6A525763", x"466E6C55", x"6C645260", x"626A4C47", x"605A5F60", x"7D8B5D6A",
									 -- x"59746558", x"645A4C54", x"5C536D52", x"515B3452", x"42585B61", x"4D506250", x"68876770", x"7D585747",
									 -- x"464C4643", x"4242445D", x"58553635", x"42383E50", x"58403E36", x"3C474658", x"5D3F4152", x"48434F51",
									 -- x"4249544C", x"3B465552", x"614E474F", x"50565257", x"605B455A", x"4C4F544E", x"51584B32", x"3D483C3C",
									 -- x"42413E4D", x"44403C2E", x"534D4343", x"3B224446", x"444A4040", x"3A3B3239", x"434C5353", x"3B4A5146",
									 -- x"4B424240", x"4C472F46", x"38444644", x"4D424841", x"404E3547", x"47523B2E", x"4039363D", x"2E423B37",
									 -- x"38423E16", x"2D412E2D", x"3E474644", x"443A384C", x"383D504C", x"54716268", x"54575D5D", x"52584A47",
									 -- x"674F3430", x"34222838", x"2A394636", x"3E493C42", x"4F55274E", x"7160724A", x"25493D28", x"464A5248",
									 -- x"5932564A", x"4147373E", x"3E434831", x"303A3D41", x"353B473A", x"4442412B", x"1F352026", x"222C4D2D",
									 -- x"13291E22", x"25322634", x"2F333032", x"37354837", x"31373B4C", x"23252F30", x"26342C28", x"352A262D",
									 -- x"2235343C", x"3233193D", x"44343034", x"29393F3A", x"31382630", x"382E4237", x"2E273632", x"43193D30",
									 -- x"373E2F3A", x"3735202A", x"35311E2C", x"251B312B", x"2127442D", x"2F2C2B2A", x"39453326", x"3236232F",
									 -- x"1E261C46", x"49313033", x"3324282F", x"2F2E4340", x"2B3F2C31", x"3C3B2739", x"33213A43", x"4E43503E",
									 -- x"3C23535A", x"375B3438", x"473C164B", x"202E3E4B", x"9560602F", x"443C4345", x"3D48472F", x"2F4B5346",
									 -- x"2A624356", x"46555E3E", x"48434049", x"3D455E53", x"3D4F4C33", x"4733435E", x"4229534F", x"4C5F4B45",
									 -- x"5750465B", x"684F4658", x"52467A47", x"4F505144", x"5D554E42", x"4E484C45", x"37355B24", x"60304B46",
									 -- x"4B51516F", x"504F653A", x"64433A4A", x"4E4B4345", x"4551442D", x"3B655A3C", x"51502C41", x"5657376D",
									 -- x"5B494D59", x"6E60715D", x"777B6154", x"42432B37", x"725D6973", x"584D816A", x"79544C6C", x"48464E57",
									 -- x"645B564E", x"4C484055", x"683B526B", x"505B4C50", x"474E6A43", x"574E4A3D", x"4443644E", x"42555160",
									 -- x"3C503D50", x"5A493B4A", x"6158665D", x"555C5974", x"815B5962", x"6D6C5D5E", x"53646050", x"655A7265",
									 -- x"5865785D", x"5C354662", x"533E4661", x"71766568", x"66666961", x"54587472", x"66605C48", x"63616269",
									 -- x"5A6A6556", x"4C4D5554", x"5450606C", x"43615569", x"5E5C696D", x"565E5951", x"706B7467", x"596A553B",
									 -- x"504A5051", x"373F5644", x"412A4242", x"20263B41", x"3D2F203A", x"47494D50", x"414A5B40", x"363D5251",
									 -- x"64455051", x"5264675D", x"604E5255", x"51535647", x"52482D45", x"51565245", x"484E313E", x"1B3A534D",
									 -- x"2D364941", x"51423F3F", x"5340373B", x"4C583446", x"3D464E37", x"3F374342", x"46434A4B", x"474C4D40",
									 -- x"3E353B2E", x"57505049", x"3D464E43", x"4B3F2F41", x"45534B3A", x"5332373F", x"3B503438", x"40404539",
									 -- x"41345835", x"403B3B44", x"34444C57", x"4B3A5346", x"4E567355", x"56551D5B", x"4B2D4F58", x"4D657245",
									 -- x"333D143A", x"4943513E", x"47513E43", x"3F413F41", x"423E4E50", x"363B4839", x"2C554752", x"6D4A3241",
									 -- x"48363D3E", x"49493B36", x"3B4A3D50", x"37373F1F", x"2F2E342C", x"272A271D", x"132F392F", x"231E240A",
									 -- x"2E24253C", x"3C342F37", x"3427252D", x"47322436", x"2D2D253B", x"3439382C", x"2C3E482A", x"1E2B3240",
									 -- x"352D253E", x"2F3B333E", x"43353E2A", x"3430343E", x"3D322A38", x"2F404A25", x"3B2D2E3C", x"31223E2A",
									 -- x"2530242E", x"492A1229", x"35371213", x"3230233B", x"33413726", x"2C331333", x"382B2F3C", x"2E2C2F27",
									 -- x"302E3543", x"3123195C", x"333E3F35", x"35402E36", x"244A2421", x"33323B60", x"44283B3F", x"405D465E",
									 -- x"26314524", x"29453A35", x"3D323639", x"322A434A", x"3B573D30", x"453C4B46", x"2A4B5237", x"3F4D4C3D",
									 -- x"4B23374C", x"2F414847", x"4E4F6942", x"435A5772", x"6F47455B", x"57646E58", x"514C4447", x"5F684448",
									 -- x"5B4D6156", x"52545760", x"585D764B", x"57535650", x"5C505145", x"4B645E42", x"47736F3A", x"3D534B43",
									 -- x"71645751", x"374E476A", x"57424740", x"515E4A45", x"4A4A5153", x"59585B4F", x"637A3C51", x"4D644F4E",
									 -- x"55425B5D", x"7261733D", x"31607554", x"416B522E", x"54645445", x"506F6D63", x"6E645B4A", x"395B4D4C",
									 -- x"556D5741", x"50655641", x"6B622C47", x"31635664", x"625D8955", x"74635B5B", x"5F514A45", x"3C645D53",
									 -- x"594E594E", x"20453A41", x"41354A65", x"6056475E", x"4C365961", x"5357494A", x"525D635A", x"5D6B6C73",
									 -- x"71606A64", x"8066647A", x"6E74686B", x"7A624964", x"5D6C6F67", x"5A3E5D7B", x"636A6F65", x"6756605C",
									 -- x"5765645D", x"534A535F", x"564F445F", x"5664776C", x"6C4D5F65", x"6B6E605E", x"60737069", x"75686D64",
									 -- x"49594442", x"4A464F40", x"3D4E604B", x"3A48443A", x"313F334F", x"5554584A", x"4D3D3035", x"484C3E3B",
									 -- x"402A384A", x"5A637462", x"6C4C565D", x"56525F3C", x"2B3A3A4E", x"554C414A", x"3B3B4156", x"37395134",
									 -- x"3F56462C", x"553E3F38", x"4C5C3844", x"40413B43", x"343D3D3B", x"3D43403A", x"463F453E", x"3E49433E",
									 -- x"473F4E53", x"393F5D3D", x"3E444547", x"4342393A", x"46334B4F", x"37425E51", x"4F41323C", x"33284C3B",
									 -- x"3D2C5241", x"4F495353", x"45445D50", x"4B575E4E", x"495D7472", x"54515253", x"4E55554E", x"4B494A23",
									 -- x"42664947", x"1F444B57", x"31524546", x"62583D27", x"32465B43", x"374A4B51", x"4750534D", x"4B39422E",
									 -- x"41363B3D", x"20212C21", x"360C263B", x"26302044", x"3136352E", x"11232329", x"1E2F2E35", x"33281F25",
									 -- x"29152E3D", x"4D2F0E45", x"31273236", x"3C39322B", x"18282B32", x"342D3238", x"35323629", x"212E2F31",
									 -- x"352B3942", x"3D395B57", x"393A3E33", x"3E373B3A", x"5F21302F", x"353E382A", x"38263727", x"2B3C3430",
									 -- x"43583F19", x"3234332A", x"2B37303D", x"2F242924", x"1E41123E", x"262E553C", x"321D1F3A", x"413B4138",
									 -- x"37292C24", x"292F374E", x"40354B46", x"1C323D29", x"374D533D", x"2C3D3C47", x"393C3433", x"44433740",
									 -- x"1E374E30", x"43433743", x"464B4A43", x"40664750", x"55595054", x"4B4A453B", x"4231283A", x"39474E52",
									 -- x"3045304F", x"4D4C5A49", x"3B5E545A", x"474E4858", x"4C4E5968", x"896C6C6F", x"7C54425B", x"6D78767A",
									 -- x"736B726A", x"6374614B", x"584F634D", x"4A3A3838", x"3C2D484C", x"31494643", x"6A538979", x"57487072",
									 -- x"41365248", x"4A514A5A", x"513A5835", x"45394D4E", x"564E4F6A", x"586D3E45", x"6E5F474C", x"623A4442",
									 -- x"39514B43", x"34575228", x"4F5B4732", x"6E66584F", x"2E2F464B", x"54484352", x"3A526F59", x"4F5A4D31",
									 -- x"475C3B45", x"504E5858", x"556E5D5C", x"52667F69", x"57585C55", x"615D6357", x"55705E47", x"485E5652",
									 -- x"60605D50", x"323F2625", x"423C484F", x"65636957", x"3F4A4F56", x"4958543F", x"4656664C", x"42565965",
									 -- x"6E44555A", x"525C5D64", x"67897273", x"6563786A", x"715E5D82", x"64616063", x"64636274", x"5A543663",
									 -- x"575B524F", x"4E464E5D", x"63647768", x"6960727D", x"796D7278", x"75758971", x"51707765", x"7865686E",
									 -- x"4F49474F", x"403E5B43", x"4F594C45", x"4B575434", x"464F4D53", x"4745494F", x"4D4A4339", x"4E484744",
									 -- x"2D474349", x"525D7E52", x"664D6453", x"4B3E3549", x"4B5A4236", x"48625644", x"3B3E5C56", x"433C474C",
									 -- x"46503B2C", x"4D3E2E38", x"4244204B", x"4E345039", x"42403E45", x"43454143", x"41302D3A", x"3E463036",
									 -- x"41463946", x"42444A3D", x"3F40374A", x"3B45542F", x"413E3A43", x"44664937", x"57373B3D", x"373D5644",
									 -- x"3D3B4242", x"5453525C", x"6C536653", x"4A6A7252", x"4F71565A", x"5A4C5656", x"505B6B56", x"465C4C4A",
									 -- x"6D604D3D", x"3A4D3C30", x"424F454D", x"536E5043", x"394E4E47", x"39436651", x"41364B5B", x"43404D39",
									 -- x"353A403A", x"31352840", x"3E323439", x"3423375C", x"2B37413F", x"1C32323C", x"363D3E54", x"26202E2C",
									 -- x"3B2D3B36", x"29231E33", x"182A2C2E", x"252B3B23", x"37312821", x"2E251F22", x"1E32292E", x"2A252E2C",
									 -- x"403F4342", x"3E334640", x"2C4E2E33", x"32333239", x"30332C5A", x"3432212F", x"3942362D", x"502A3732",
									 -- x"353D393B", x"39364447", x"41494D4D", x"363A3431", x"2A281C22", x"173C320E", x"16321F13", x"35282C33",
									 -- x"33374D50", x"31323825", x"3C3C383A", x"3A31443A", x"535C4E3A", x"4159462D", x"283F292A", x"3E354338",
									 -- x"426B323E", x"584B5B4F", x"644A2D40", x"314B4A2E", x"5F505759", x"4C4C5651", x"4C693D45", x"4F64414E",
									 -- x"48555B65", x"644E443A", x"30594B4A", x"426D5B2D", x"544F5D5D", x"6D4D5D61", x"74606460", x"5F534753",
									 -- x"5660435F", x"50504E5A", x"42516A38", x"42483F42", x"53585A6D", x"43845837", x"615A6E37", x"5A5C6B5A",
									 -- x"6652534F", x"454A6746", x"40225960", x"5337545A", x"58473F49", x"41424C67", x"554B3260", x"64604349",
									 -- x"4959503F", x"3986434C", x"574C384A", x"57527E5D", x"584B544D", x"7B364459", x"504F584F", x"4F65425B",
									 -- x"553E584D", x"56703344", x"38554E73", x"6F5F7F6E", x"5C464D53", x"3A4F7659", x"486B645F", x"4B5E4654",
									 -- x"655C5546", x"54453853", x"37353B4D", x"4B3F4F50", x"4D564B4E", x"4D4E3950", x"4C544F5F", x"54564A47",
									 -- x"6A4E4958", x"5C3F614D", x"60655C6D", x"5A5E6B64", x"5D5B5553", x"4B634F4D", x"655E6082", x"6A594052",
									 -- x"5B605354", x"63666667", x"70647381", x"61767063", x"62727579", x"787A8682", x"7781976D", x"6B836C71",
									 -- x"534E4D41", x"38394A45", x"46543E40", x"574D4852", x"514E5052", x"47434351", x"50434E5A", x"6C4B534F",
									 -- x"4E69504E", x"5164693E", x"2F350F43", x"5740644E", x"4E4F4B3C", x"47354837", x"2C383D50", x"435B404D",
									 -- x"27364547", x"4343404E", x"3B223D41", x"3D363643", x"352E3531", x"38313B3B", x"4A383049", x"59514144",
									 -- x"3C3B403F", x"3C3C4240", x"422C3D39", x"3040352D", x"4D424528", x"4C4B402D", x"32353639", x"4751463A",
									 -- x"3F3A474D", x"4A4C5352", x"46404D57", x"586E805B", x"56694C30", x"30484F47", x"34425945", x"4C68465C",
									 -- x"4451425F", x"5C454A35", x"583E4A85", x"3C4D474B", x"403E3A2D", x"4041444F", x"353B4749", x"363C404D",
									 -- x"38415747", x"444C3132", x"3A3A4237", x"44444541", x"412F3B3B", x"2E32353C", x"4E1E3430", x"1336372C",
									 -- x"17253730", x"242B3A1B", x"21310F24", x"3E2D203A", x"352C3633", x"2F2A2128", x"363D1F20", x"242D372E",
									 -- x"3E352D30", x"2B342421", x"374E3730", x"3139313E", x"355A3E47", x"32384B2E", x"35363635", x"36381D41",
									 -- x"2C453B37", x"31384649", x"34263338", x"294A473F", x"4C274037", x"1E2D2D29", x"4F4F3C34", x"5A45411E",
									 -- x"2B432E5F", x"47395232", x"3B342D3A", x"3F2B3930", x"2E3F3C2D", x"674F453A", x"3A485060", x"445E4835",
									 -- x"59453F65", x"2B284C5A", x"2B423F58", x"534B5C38", x"635C2968", x"654B5242", x"514F5154", x"4E505B4F",
									 -- x"5A674E48", x"5C585449", x"49664D56", x"785F6563", x"636D6870", x"595C495E", x"605F5D5A", x"71785552",
									 -- x"415E627C", x"43394E43", x"4460655D", x"4B504674", x"5C505F70", x"5C453F48", x"4D53755C", x"42484029",
									 -- x"545C644E", x"58583747", x"5C577062", x"3F5B6C5D", x"5F563B5B", x"5D5D654C", x"54451773", x"65475E59",
									 -- x"60596762", x"5A873D62", x"583F375A", x"65527D6D", x"4A646056", x"543E6272", x"38576E4E", x"3A593268",
									 -- x"4E3D5C4F", x"3445366D", x"65346834", x"472F2A5E", x"44545652", x"4B50573E", x"59804B5C", x"4C675A3F",
									 -- x"5F2D5254", x"5452544E", x"40474528", x"38566C48", x"34585E3F", x"53714444", x"4D335853", x"7355422F",
									 -- x"52594C5B", x"74466F59", x"705F575E", x"5E5C4A69", x"543F5E48", x"3A4D4038", x"64605D68", x"75666B49",
									 -- x"56766769", x"91886C71", x"6669658A", x"5974785B", x"5B696D66", x"71626170", x"91B0907A", x"86938B89",
									 -- x"5152492A", x"40534C51", x"554C5152", x"544C3A40", x"5C594840", x"40454940", x"5252526B", x"5B525340",
									 -- x"464C4755", x"41443043", x"41294364", x"33425A44", x"4B523641", x"35404A20", x"37424F42", x"463E4845",
									 -- x"415D595B", x"46495E26", x"30405340", x"3E3D3837", x"2D282A23", x"2A2A2818", x"32353031", x"4839423A",
									 -- x"312F2D26", x"2C3C292E", x"2F273030", x"3C302940", x"39372C26", x"3D40363E", x"253A222F", x"3635313A",
									 -- x"102C3724", x"3C3A3437", x"34483F3F", x"504E4A4B", x"4742434C", x"45494C55", x"4F453F3D", x"3D3C4626",
									 -- x"45476750", x"413A2C31", x"1C372A59", x"4345393E", x"45392F30", x"3F263143", x"2C2E391D", x"373A352E",
									 -- x"33363D30", x"331A0F37", x"4F303B37", x"2C373234", x"4C162630", x"422D2C2E", x"371D3129", x"3B2D2C2B",
									 -- x"26324C2C", x"33282422", x"25211D2A", x"232E2735", x"2B1A3038", x"2B35303A", x"3A2F2827", x"1D2F3A3F",
									 -- x"351C2C25", x"24342A2B", x"3C19422F", x"40595649", x"3F383C49", x"42524B26", x"1A413D4F", x"36373D2C",
									 -- x"29513420", x"3C433C36", x"1B3E2E3E", x"403C3630", x"413A452F", x"3435252A", x"3D38353F", x"5A1E3141",
									 -- x"31353133", x"3D3A3C4C", x"473F4955", x"3F3B3E45", x"3C394344", x"5A4B3366", x"53554A53", x"433C8A4B",
									 -- x"593E495A", x"243D3E37", x"4E4A6861", x"5C57615F", x"6B535160", x"63545052", x"4F685346", x"49545B64",
									 -- x"544C4176", x"575A5655", x"545C6B51", x"645C626C", x"73738E7A", x"776D5856", x"6C7F6F6A", x"50595C7B",
									 -- x"61635758", x"5E656A51", x"5D6B6D71", x"5E586863", x"5A5D4E52", x"4C37414F", x"5440605A", x"5C434763",
									 -- x"56504E2F", x"5D482443", x"4B415A59", x"484A474F", x"6A5C6967", x"6254664E", x"49676376", x"3942814B",
									 -- x"37747E74", x"39595751", x"46505162", x"54453D53", x"72735863", x"7A4D3D5A", x"504B5A40", x"45454440",
									 -- x"5E677863", x"44636271", x"554A7051", x"64394D51", x"30683044", x"4D53502C", x"5C7B503A", x"47574E5D",
									 -- x"63576D65", x"5C57554D", x"46434D4A", x"4B5E5E4E", x"5C605857", x"614E3B45", x"58636255", x"5B4F6B58",
									 -- x"51535555", x"516B624E", x"556A5A4D", x"54584E52", x"5C435F51", x"57835C4F", x"4B656D56", x"72746E71",
									 -- x"6E726E74", x"7A767067", x"6E796E67", x"77707261", x"525A5C58", x"6347796A", x"7978656A", x"6F768678",
									 -- x"4C4F3943", x"49494B49", x"5457504D", x"5260514A", x"552A3A4E", x"3E324740", x"4C545945", x"433F5653",
									 -- x"4B564C52", x"52342A3E", x"323F6C48", x"48474E51", x"46474C32", x"4757574E", x"54486641", x"304A4C4F",
									 -- x"564C443C", x"443B3E31", x"33403B3B", x"362A2218", x"2D292336", x"29293634", x"3A4D3626", x"67384635",
									 -- x"352B312E", x"32272326", x"2C333527", x"3B2D3139", x"314E364E", x"58374242", x"353D223B", x"49310F36",
									 -- x"2F3D3734", x"3D2B342C", x"3D233C3F", x"434E3E44", x"403D3A43", x"403A423D", x"404A3B24", x"48463122",
									 -- x"383E4744", x"2D41292C", x"3048553A", x"32474332", x"373C2A37", x"48454036", x"272F2927", x"36351E1A",
									 -- x"36463437", x"351E2428", x"412D2F2D", x"27372D40", x"4F4F1D32", x"57143929", x"2A411631", x"332B2634",
									 -- x"36312D38", x"382B3B27", x"2E262B21", x"241F0E1F", x"290F282C", x"302A353B", x"29241D20", x"2B283434",
									 -- x"32213A34", x"313B3E34", x"35332E2F", x"373C3337", x"2C403238", x"44414A51", x"73434B46", x"4D34465A",
									 -- x"3847463F", x"5B4C443B", x"26393154", x"3E1E4136", x"322C3836", x"3B342D42", x"182D342E", x"0F313329",
									 -- x"2A313221", x"3334304A", x"5843392E", x"55595559", x"62523868", x"4B4B5556", x"78685945", x"456A5149",
									 -- x"5C4F626A", x"4651463D", x"535E544C", x"4B4E5761", x"4B515554", x"59565C55", x"3A6E514B", x"4B675563",
									 -- x"5B4F4958", x"4F474E34", x"4465474D", x"5659686C", x"6D605A63", x"7F72615C", x"5A75693D", x"5139343A",
									 -- x"5A5E6860", x"4D576F71", x"5F6B5A5F", x"79666857", x"55512F4F", x"403A5D5B", x"56615755", x"56554348",
									 -- x"43433E38", x"42514743", x"4C38484C", x"4A493A3C", x"4C45724E", x"42393141", x"394A5D6C", x"536C3742",
									 -- x"51585750", x"55614E25", x"4E4D5A63", x"4D4B464F", x"3055504A", x"4A566A43", x"474D4650", x"3062555D",
									 -- x"665F6D3C", x"52605857", x"4E3C5C61", x"777C6B41", x"445D6431", x"53526C61", x"79765E4B", x"845D7864",
									 -- x"51747F68", x"54676E4F", x"464A5260", x"52455468", x"5361666B", x"5068534C", x"4F6D494E", x"494C605A",
									 -- x"42545855", x"5F5B5356", x"42535E64", x"5D5F5662", x"66597354", x"59696955", x"57537765", x"6862715C",
									 -- x"6261574A", x"535C6262", x"775E5263", x"53426A4A", x"47513D3C", x"5B546658", x"5D575F4F", x"5C776973",
									 -- x"564D5055", x"4F5C5441", x"494D564E", x"3F4A4F4E", x"46405036", x"3F4B3B4D", x"31534F40", x"3349544E",
									 -- x"473E4651", x"48283B47", x"26363D55", x"4F414348", x"2A48494D", x"53495561", x"32476E3C", x"4E3B433E",
									 -- x"44402E3E", x"2D2A1E4D", x"45432755", x"3636272F", x"361C363A", x"3D323F55", x"584A5939", x"37454B3C",
									 -- x"22233032", x"2A283A47", x"3C413833", x"3B343F34", x"353C4137", x"41384F40", x"42323445", x"3B28303C",
									 -- x"583F2334", x"3F343229", x"47485348", x"3B39462E", x"39302C40", x"32322132", x"290F3542", x"3E403733",
									 -- x"413F3A35", x"3837333F", x"4A404222", x"42373A3E", x"3336403E", x"46414130", x"2E223A22", x"32592937",
									 -- x"35284A33", x"161E172A", x"2E2A2331", x"2B222A30", x"4C383735", x"2E3A5B37", x"31433647", x"54372B34",
									 -- x"2328402D", x"303B2425", x"1F351C28", x"2F232A2C", x"3329272B", x"323C393D", x"3D35282B", x"33483F33",
									 -- x"33382E2C", x"3D2F3B37", x"3853442E", x"3033311A", x"30272F32", x"314A7275", x"81444849", x"613F5840",
									 -- x"2066474C", x"4E335A40", x"42333F58", x"233F272A", x"481A2E27", x"2C3C2D39", x"35252315", x"39371E2C",
									 -- x"2D3D4330", x"4F414A40", x"4B3D4C47", x"6F5E4964", x"52375133", x"3E4C5547", x"54574B52", x"454E292A",
									 -- x"4B633944", x"593B2836", x"4D5A3831", x"47525442", x"55513F3A", x"503F403D", x"4E565156", x"5D556046",
									 -- x"563A5C4F", x"4554444A", x"575F4848", x"50596973", x"605A634F", x"53554959", x"6D3E4B6F", x"60687256",
									 -- x"66766441", x"6E4F3356", x"4A535B51", x"3C505B6A", x"534A575C", x"55596E5C", x"3D595551", x"6B483B49",
									 -- x"51353D4F", x"59637551", x"5450574A", x"38403931", x"4F423F6E", x"59472F42", x"33575A42", x"544E334D",
									 -- x"39583953", x"6570344F", x"6C565950", x"5A795960", x"565A5453", x"5664545F", x"5D655F5B", x"4F565B5C",
									 -- x"4B692F56", x"72594A60", x"774D5061", x"4351685B", x"68859867", x"80698062", x"60404D49", x"5551486E",
									 -- x"54535F5F", x"57606B6F", x"565F6360", x"5A565745", x"49715D5C", x"6D6C5054", x"4D686069", x"66827847",
									 -- x"5D523E61", x"5B686166", x"775E8869", x"626A7C6D", x"67703C65", x"6F595D63", x"5156705E", x"52676351",
									 -- x"5E405135", x"42634B49", x"3B71355C", x"4943473D", x"6B567151", x"46736345", x"5B575B5F", x"687D675F",
									 -- x"4F435657", x"4F61514A", x"564B5953", x"444E5B50", x"3C473E46", x"51424D4E", x"5150545B", x"5B5C5D56",
									 -- x"594B3B5B", x"62493037", x"494D4656", x"4F573C42", x"46474B4D", x"41472E23", x"3D534A2C", x"50493F29",
									 -- x"384B444C", x"2E554249", x"2D2C432E", x"4058392F", x"51373138", x"44424E4C", x"3F1F4351", x"263B351E",
									 -- x"482A424D", x"33322F2D", x"16493B45", x"2D3B4039", x"5B223848", x"29253B32", x"37444B3E", x"3A282D1E",
									 -- x"3F3E4042", x"394A3A58", x"534F4D40", x"3D364234", x"2B361838", x"52452232", x"1529423C", x"40503F3C",
									 -- x"484E4047", x"42372D33", x"3E4B4236", x"34323846", x"1C274F4A", x"3F3F382A", x"3F29482D", x"2C372F40",
									 -- x"2B232329", x"1919302A", x"411E2627", x"281D2E35", x"22303037", x"26383A04", x"2E31423E", x"38353529",
									 -- x"25565330", x"28313032", x"302B2D3F", x"383E5033", x"3A2E103B", x"4231283E", x"3E5C3729", x"362F3052",
									 -- x"4314231D", x"3D203424", x"23303125", x"2F351933", x"49394237", x"363F4638", x"26341E1C", x"3F4E3E3C",
									 -- x"3E284537", x"4A4F4F3E", x"3C5C456A", x"2A51342F", x"39383026", x"233B2F32", x"260E323A", x"36493B39",
									 -- x"523D423F", x"37454947", x"65475971", x"6D513B5B", x"2643674D", x"473D3B4B", x"4B3F1F70", x"453D3A3B",
									 -- x"53474F4F", x"455C4843", x"4F505845", x"325B4531", x"4D44393C", x"56483847", x"51416E4F", x"6B374643",
									 -- x"414A4E4A", x"74545543", x"4E59544A", x"4A5D4D61", x"69574A41", x"61635770", x"4B5C799C", x"645C5A6B",
									 -- x"57636551", x"5E5A3B44", x"605C45B5", x"A76D4459", x"52645659", x"67634F65", x"5866605B", x"564C4861",
									 -- x"4A5D4A39", x"5B5B4E54", x"6E58645D", x"4D714F51", x"4F4D4B44", x"5E526E6E", x"5B6F5C62", x"635B6862",
									 -- x"4B4B6A6F", x"5C563D6D", x"56586762", x"5C407163", x"6F70737E", x"61525568", x"687B5E4A", x"4C385672",
									 -- x"57716153", x"4E724455", x"34444863", x"59535861", x"456D5E54", x"61575D65", x"3E535B49", x"42534936",
									 -- x"5A5D657C", x"6C64655C", x"4D645D59", x"76596055", x"62777286", x"96827A6E", x"71987AA5", x"7C7B736E",
									 -- x"606D6261", x"6466645F", x"824A6D71", x"59586359", x"5F806372", x"79626074", x"504D6132", x"554D4949",
									 -- x"5C26464C", x"1652594D", x"47434921", x"4A655E55", x"62636F79", x"50525F56", x"46664166", x"78426170",
									 -- x"41435759", x"54523B4E", x"63464A52", x"6166542B", x"44443653", x"6A534E50", x"52715E60", x"82623E44",
									 -- x"5B4C524D", x"2D475758", x"514D4457", x"523C2A39", x"3644432E", x"28351D37", x"464D5066", x"59524E46",
									 -- x"3C476338", x"40453435", x"45503C23", x"30423A3F", x"463C4149", x"4D313A35", x"40394041", x"2E443B45",
									 -- x"5B294545", x"27443D34", x"2F522D37", x"2B3D3131", x"4E34272A", x"3E3D372E", x"3D543239", x"3D543423",
									 -- x"24404858", x"5C3B4166", x"4455323A", x"463B554C", x"27244946", x"40332632", x"3B3E4935", x"4151373B",
									 -- x"40523A38", x"37362C3D", x"3F2E3A37", x"32303733", x"17344F29", x"072E271E", x"613E1F1E", x"3A2C2030",
									 -- x"33291F1A", x"23242236", x"2C342819", x"294C3B39", x"3D3D362D", x"314A2C29", x"44424C34", x"22333133",
									 -- x"30513C2C", x"2A2B2A32", x"3D434940", x"44413D2D", x"3153322B", x"262E3E37", x"34403345", x"43233F16",
									 -- x"38182B32", x"57372A1F", x"26112328", x"2B51344B", x"4F36322E", x"3A2F3638", x"51383F27", x"5151464A",
									 -- x"42524E25", x"4D314B48", x"4019333E", x"3455332C", x"3B3E253D", x"3C473A48", x"3B4C5731", x"38363C47",
									 -- x"4F604715", x"444F403F", x"56464F4C", x"4935383E", x"4B565F49", x"45516E5A", x"4C375468", x"254B594C",
									 -- x"4F7B574B", x"4A4F3944", x"4C433150", x"38525857", x"34364B43", x"44685E5D", x"6F4E5C57", x"524D5868",
									 -- x"626C3D4D", x"5C5C5D55", x"5D5D566E", x"535A6372", x"7E76605E", x"72565D69", x"6B786D5B", x"294A575E",
									 -- x"50627476", x"615F5C73", x"6364657A", x"9D7D5C4C", x"55533C4D", x"55584150", x"7A5D5952", x"3F5A585A",
									 -- x"59696751", x"59715670", x"6646586B", x"6F5C5158", x"464A554A", x"6E4E4D7B", x"5C70554E", x"60436544",
									 -- x"62683A58", x"4240735B", x"2E4A6260", x"5A4A5D41", x"53725C65", x"4B535B5C", x"5956364F", x"4639455B",
									 -- x"684F6650", x"46585370", x"6A6F6681", x"64555265", x"47363E3C", x"5A645060", x"5C6B4333", x"8E794C6D",
									 -- x"6B7D6A64", x"9C6E5E60", x"515F4B63", x"6E687766", x"73968497", x"945D6F70", x"684E5577", x"6E5C6664",
									 -- x"8D5B6869", x"56415A59", x"5155507C", x"5E424E38", x"3E3B3052", x"6C4A5656", x"4B4D4B48", x"47413756",
									 -- x"51514553", x"6C534436", x"7B555663", x"515D4D58", x"60645B72", x"5A384379", x"52627647", x"67605C7B",
									 -- x"4A4F5454", x"4C4C485E", x"61555446", x"47464949", x"3F455262", x"575C7060", x"4D684858", x"4E414353",
									 -- x"57305345", x"4C474E5F", x"54474F47", x"44453C64", x"42373139", x"38393732", x"48635435", x"4A4E403C",
									 -- x"44443352", x"37415B3B", x"4342202D", x"2736435C", x"39305627", x"392C3A38", x"323E643D", x"1E3B3834",
									 -- x"1016393F", x"31483D2D", x"433A2938", x"3D38241C", x"30463919", x"47374E3D", x"472F3B47", x"50383322",
									 -- x"353E483E", x"42454A64", x"503E3A47", x"342A2244", x"54414441", x"39132F36", x"3A363F1C", x"4259363E",
									 -- x"3A354545", x"1B2B4248", x"3734274D", x"430E4534", x"26334426", x"0E2C344D", x"49373D3A", x"32442C32",
									 -- x"3C3E4A2E", x"333D2A55", x"46322A31", x"423F4F40", x"40342F25", x"273B3534", x"33413D24", x"37382957",
									 -- x"37341940", x"543E3433", x"21484133", x"35413F36", x"503A332E", x"4C594D37", x"2D3E4E5F", x"43296338",
									 -- x"3F372251", x"3A38353C", x"3F41372B", x"34362E41", x"452F3349", x"52353C32", x"42404862", x"5C603442",
									 -- x"4A623B6C", x"495B2647", x"47624D4C", x"41373A44", x"44354235", x"3848443A", x"433C3739", x"363D5C3E",
									 -- x"35715F4E", x"6744472F", x"3C484B45", x"47361529", x"4257574E", x"4649505D", x"3E3F7B64", x"4A47544D",
									 -- x"587E5145", x"4B414450", x"40644145", x"484C4C45", x"3557564B", x"6D664A5A", x"36464557", x"694C5C56",
									 -- x"595D5068", x"46486B51", x"4A656E56", x"576B545F", x"66657171", x"6143583D", x"5A535F5E", x"5B807F59",
									 -- x"66806B6A", x"8C583F69", x"6E62684B", x"4336505F", x"4C465959", x"6F735554", x"64506E5F", x"594C6456",
									 -- x"544F675E", x"47514D6B", x"67637D6C", x"59725F77", x"5948584F", x"3B545250", x"4B494E43", x"4C586B3B",
									 -- x"6753607A", x"63564F4E", x"4B3B7272", x"785C8B46", x"3C3C6155", x"60466E5F", x"62584472", x"3C595B64",
									 -- x"5D5F6B5E", x"756E5849", x"585B8369", x"6041686D", x"602E5649", x"40746E66", x"65564E58", x"78727474",
									 -- x"72667B62", x"5470815E", x"54595C59", x"775E657F", x"767E8060", x"64655764", x"546E5851", x"5331534D",
									 -- x"595E6854", x"32565F63", x"64545E57", x"462F4464", x"51302F54", x"6D515F5D", x"60432856", x"3654564C",
									 -- x"45625657", x"69595649", x"58523E56", x"5F5E543A", x"465D5557", x"59515458", x"4E577948", x"55656D59",
									 -- x"5D595554", x"46545F58", x"5B554F47", x"504F4A52", x"4E706055", x"55555959", x"53226C69", x"35534C54",
									 -- x"49477142", x"4149454A", x"2D4A354B", x"4B484C3D", x"33414B3E", x"4D4A3A43", x"582E282E", x"414C4F48",
									 -- x"452E4133", x"45514936", x"38212A38", x"4240422C", x"3735472C", x"3E414032", x"1340482B", x"41383959",
									 -- x"3B483543", x"4F43413E", x"3A302A39", x"23363736", x"3C484134", x"2D18453D", x"36434C43", x"1E4E4F3F",
									 -- x"414A4827", x"37457857", x"31232B55", x"383C4052", x"36423B1E", x"323C3532", x"433D2D36", x"5F464047",
									 -- x"36402941", x"374A2940", x"4E3E3A28", x"28314047", x"3A314431", x"2E253753", x"2A255B4F", x"341C2A4F",
									 -- x"293A3A32", x"323A4240", x"4D2C3C36", x"3B37463D", x"2438372E", x"2B2B3D1C", x"283B3B1C", x"372A2143",
									 -- x"34183E39", x"43502042", x"46342F47", x"3B45294C", x"3E1A483B", x"596E483E", x"2A614814", x"18283530",
									 -- x"3B45455B", x"29504434", x"45454122", x"483D4044", x"2045493E", x"3D314648", x"3D394547", x"45314434",
									 -- x"47494B5C", x"325D4741", x"42513347", x"37393F2F", x"524B3C56", x"3F402D36", x"4339162D", x"20354A31",
									 -- x"55442141", x"5B4E4D36", x"35344E41", x"45462B41", x"4C4B4661", x"4F43494F", x"4A5E362D", x"5C544F4A",
									 -- x"6F153B47", x"37374C65", x"3A505F62", x"6E37303D", x"3D453F49", x"613B4326", x"5439294F", x"5163693C",
									 -- x"5C4F497E", x"57835330", x"624D4E34", x"54453F64", x"6763483F", x"5B59565F", x"5F536760", x"665B6068",
									 -- x"5D644C4B", x"54595D4D", x"4F53545C", x"526B4245", x"434F4661", x"50466C5A", x"5C7E4775", x"74774A55",
									 -- x"5A4D5B4D", x"403A5650", x"576F614E", x"425D5750", x"645E5455", x"60594D4F", x"4A3C665E", x"4461474A",
									 -- x"5E4D5863", x"7467525D", x"4B497C7C", x"786B663C", x"817D525A", x"656E8067", x"6E647B71", x"6F4F677C",
									 -- x"4357645C", x"62726678", x"614C7D5A", x"6C416850", x"415A6169", x"476A7E46", x"576F515A", x"564E4C85",
									 -- x"655C445F", x"51326B71", x"5F497457", x"5C5A5962", x"6F6A4950", x"654A5852", x"645E6159", x"40525653",
									 -- x"3667655B", x"55674D78", x"6860505E", x"511F5665", x"555A755B", x"613E5B64", x"44414A59", x"49496D51",
									 -- x"45555C74", x"5C562C52", x"574E434C", x"575D4F52", x"533E6B6C", x"5A605A57", x"594C6064", x"6C736E6C",
									 -- x"5F5E6062", x"555D533A", x"58564F49", x"494C4F63", x"5D504A5C", x"67675455", x"4F526555", x"4D4C6148",
									 -- x"38515F42", x"484E3A53", x"4E4E3E56", x"504F4440", x"45465D38", x"36514347", x"31303C52", x"43413841",
									 -- x"2E244444", x"433D4741", x"3F372149", x"56424827", x"4C49374B", x"3C3E3A4E", x"384D3C3D", x"5036404A",
									 -- x"684F3246", x"533C4140", x"38403442", x"36403E3C", x"464B2F32", x"2A373334", x"473E4842", x"33473237",
									 -- x"4B483B52", x"3D644549", x"4D4C5646", x"35644336", x"37312E42", x"26235B66", x"4840303E", x"3C2B3F1B",
									 -- x"2E433345", x"2937334D", x"3C4F7049", x"3E414D3D", x"363E4E31", x"363B5845", x"20463F0D", x"35263537",
									 -- x"34323531", x"2D383929", x"28242B3D", x"3B49164B", x"2C3B4C29", x"2C3D473B", x"2B3D4532", x"38384140",
									 -- x"313F5638", x"333B2B40", x"3C424136", x"496D324F", x"6644583E", x"3A441E22", x"33343737", x"3E303047",
									 -- x"46384040", x"3B391848", x"43406945", x"39375940", x"385E4D34", x"4B595344", x"3D3D3927", x"602B4440",
									 -- x"513B4142", x"4858323C", x"6545414B", x"623F4141", x"41443830", x"5A374326", x"3B3D3D34", x"382D302F",
									 -- x"521F3A47", x"57566642", x"5F496237", x"404A674E", x"2B4A553A", x"5E424447", x"4D5F4C5E", x"654B336A",
									 -- x"524D4D31", x"3A484C53", x"4D595353", x"63324D3A", x"36514131", x"45495F34", x"6147503B", x"514E5B57",
									 -- x"5F78586E", x"5658584D", x"775D566C", x"6D529068", x"6C614F66", x"59615F59", x"573F5E62", x"5F4B4F55",
									 -- x"514C6774", x"2D516C2F", x"346B555D", x"614F4B32", x"434D555B", x"525A374B", x"56514558", x"49514F31",
									 -- x"57634A30", x"6867695E", x"403A5340", x"6F5C5756", x"585B4755", x"614E4146", x"6C1E5859", x"55745F3F",
									 -- x"587F5647", x"5F66596D", x"5C556558", x"7481A361", x"72B26F54", x"73736F59", x"456D5430", x"3157504A",
									 -- x"5A544746", x"4A58533E", x"5F35465D", x"33286578", x"52795549", x"5647743E", x"453F5150", x"445D3E60",
									 -- x"56506556", x"9D675E6E", x"616B6452", x"4474553C", x"6492834A", x"64565242", x"5942645D", x"59585E63",
									 -- x"70695A62", x"6E635660", x"5C716260", x"51446161", x"4E616755", x"591E5656", x"354B5D6D", x"7257625C",
									 -- x"455A594A", x"5D78553D", x"577A7F70", x"5A55727B", x"62747F6B", x"4D587858", x"60574D5B", x"71806F72",
									 -- x"5B5C585A", x"5E634F4B", x"5A5A5A58", x"4A4C4D60", x"51604987", x"7E445452", x"525A504F", x"5B545264",
									 -- x"41325651", x"454F695A", x"454E4C45", x"363B3D3D", x"3A46493A", x"44534C4D", x"48493C49", x"473D3546",
									 -- x"3450433A", x"432A4C3C", x"41503B33", x"46464146", x"41505449", x"35573D46", x"4E504B32", x"2A47482D",
									 -- x"43223E4B", x"3B394536", x"42483830", x"5724354A", x"4F323643", x"32473A3D", x"473E5C45", x"3A433741",
									 -- x"42454E3B", x"523E2E47", x"3C413227", x"39583742", x"3B333848", x"353B5935", x"54393938", x"41402A3F",
									 -- x"4F434B3E", x"372E5A3A", x"43453F63", x"30333D2B", x"37394948", x"40384922", x"2F332C39", x"423F4034",
									 -- x"34353A3A", x"2B242D33", x"30264237", x"31424239", x"2E394941", x"4040533B", x"364C494E", x"45434545",
									 -- x"3754483B", x"4736332C", x"393A494B", x"53503A3C", x"444A4948", x"3136354F", x"37263E41", x"3F375843",
									 -- x"354D523D", x"2F382A3C", x"3E37233F", x"5B374030", x"37414B42", x"373B3B3B", x"3C4D4E36", x"3C384638",
									 -- x"63443740", x"4C5D3C40", x"554C4D54", x"33404949", x"4D414745", x"4E465249", x"4D44514D", x"46483C63",
									 -- x"4D555154", x"5D363154", x"574B2F64", x"4E50584C", x"39486933", x"47472252", x"5453515B", x"57495449",
									 -- x"46725653", x"4F4B5059", x"63635036", x"504F5A64", x"435F5B52", x"4E595049", x"4A586657", x"6245586A",
									 -- x"3C605C5E", x"3A434E65", x"65585758", x"58576657", x"41784459", x"50534958", x"4C4D5F4F", x"4D4B4A55",
									 -- x"79505463", x"4F4E5F5D", x"7254314B", x"5B515048", x"6F605455", x"60706432", x"56646345", x"57705550",
									 -- x"5B546255", x"5E696F5C", x"48756D4E", x"56636560", x"58606560", x"806A605A", x"664C564C", x"4B726453",
									 -- x"6F4D645A", x"62456182", x"5A3F5F54", x"615D556B", x"5B546068", x"6D5A5F57", x"4D504F54", x"51595641",
									 -- x"4C34443E", x"5A585A4B", x"60605452", x"62506B5E", x"696F6752", x"4D4A6078", x"5D5F6051", x"64595561",
									 -- x"59635555", x"6762826B", x"625D5B64", x"5B4F755D", x"6B5E8C4F", x"5A5F5543", x"6B3F7D5C", x"3760606B",
									 -- x"746B4A56", x"6D636157", x"3F627363", x"5C4A4B62", x"74676A5E", x"51506165", x"504B5869", x"69455C7F",
									 -- x"5577595C", x"555D705C", x"696E5667", x"6F6B6B78", x"646E695E", x"615D5760", x"60605B5C", x"585D6A69"
									-- );

	type States is(T1, T2, T3);
	signal 	RxState, TxState : States;--, MCUWrState, MCURdState

	signal	FrameRate			: std_logic_vector(31 downto 0);
	
	signal	TPGData				: std_logic_vector(31 downto 0);
	signal	NextTPGData			: std_logic;
	
	-- signal	RowCounter			: std_logic_vector(11 downto 0);
	-- signal	ColumnCounter		: std_logic_vector(11 downto 0);
	-- signal	PixelNumberCount	: std_logic_vector(31 downto 0);

BEGIN

	Avalon_Proc : process(nReset, Clk)
		begin	
			if (nReset = '0')then
				-- s0_readdatavalid <= '0';
				NextTPGData <= '0';
				s0_readdata	<= (others => '0');
			else
				if rising_edge (Clk)then
					if (s0_read = '1' and s0_chipselect = '1') then
						if (s0_address <= "00") then
							NextTPGData <= '0';
							s0_readdata <= TPGData(15 downto 0);
						else
							NextTPGData <= '1';
							s0_readdata <= TPGData(31 downto 16);
						end if;
					else
						NextTPGData <= '0';
						s0_readdata <= x"0000";
					end if;
				end if;
			end if;
		end process Avalon_Proc;

	FrameRateGenerator_Proc : process(nReset, Clk)
		begin
			if (nReset = '0') then
				FrameRate <= (others => '0');
				Int <= '0';
			else
				if rising_edge(Clk) then
					if (FrameRate = x"004C4B3F") then--25FPS
						FrameRate <= (others => '0');
						Int <= '1';
					else
						FrameRate <= FrameRate + 1;
						Int <= '0';
					end if;
				end if;
			end if;
		end process FrameRateGenerator_Proc;

	TPG_Proc : process(nReset, Clk)
		begin
			if (nReset = '0') then
				TPGData <= (others => '0');
				-- RowCounter <= (others => '0');
				-- ColumnCounter <= (others => '0');
				-- PixelNumberCount <= (others => '0');
			else
				if rising_edge(Clk) then
					-- TPGData <= VideoData(conv_integer(PixelNumberCount));
					if (Int = '1') then
						-- TPGData <= x"03020100";
						-- RowCounter <= (others => '0');
						-- ColumnCounter <= (others => '0');
						TPGData <= (others => '0');
					else
						if (NextTPGData = '1') then
							if (TPGData = (PixelNumber - 1)) then
								TPGData <= TPGData;
							else
								TPGData <= TPGData + 1;
							end if;
						else
							TPGData <= TPGData;
						end if;
						-- if (NextTPGData = '1') then
							-- if (RowCounter = (Row - 1)) then
								-- if (ColumnCounter = (Column - 1)) then
									-- TPGData <= x"00000000";
									-- RowCounter <= (Row - 1);
									-- ColumnCounter <= (Column - 1);
								-- else
									-- TPGData <= x"03020100";
									-- RowCounter <= (others => '0');
									-- ColumnCounter <= ColumnCounter + 1;
								-- end if;
							-- else
								-- TPGData(7 downto 0) <= TPGData(31 downto 24) + 1;
								-- TPGData(15 downto 8) <= TPGData(31 downto 24) + 2;
								-- TPGData(23 downto 16) <= TPGData(31 downto 24) + 3;
								-- TPGData(31 downto 24) <= TPGData(31 downto 24) + 4;
								-- RowCounter <= RowCounter + 1;
								-- ColumnCounter <= ColumnCounter;
							-- end if;
						-- end if;
					end if;
				end if;
			end if;
		end process TPG_Proc;

END Arc_TPG;

