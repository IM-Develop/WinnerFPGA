`timescale 100 ps/100 ps
(* black_box_pad_pin="REFCLKP,REFCLKN" *)module EXTREFB (
  REFCLKP,
  REFCLKN,
  REFCLKO
)
;
input REFCLKP ;
input REFCLKN ;
output REFCLKO ;
endmodule /* EXTREFB */

